`timescale 1ns / 1ps
`default_nettype none

module fsqrt_d(
  input wire [31:0] x,
  output wire [31:0] y,
  input wire clk);

  wire [0:0] swire;
  wire [7:0] ewire;
  wire [22:0] m;

  
  function [22:0] tab (
    input [11:0] M
  );
  begin
  case(M)
12'd0 : tab = 23'b01111111111101000000010;
12'd1 : tab = 23'b01111111110111000000011;
12'd2 : tab = 23'b01111111110001000001000;
12'd3 : tab = 23'b01111111101011000001110;
12'd4 : tab = 23'b01111111100101000011000;
12'd5 : tab = 23'b01111111011111000100010;
12'd6 : tab = 23'b01111111011001000110000;
12'd7 : tab = 23'b01111111010011000111111;
12'd8 : tab = 23'b01111111001101001010010;
12'd9 : tab = 23'b01111111000111001100110;
12'd10 : tab = 23'b01111111000001001111100;
12'd11 : tab = 23'b01111110111011010010100;
12'd12 : tab = 23'b01111110110101010110000;
12'd13 : tab = 23'b01111110101111011001100;
12'd14 : tab = 23'b01111110101001011101100;
12'd15 : tab = 23'b01111110100011100001100;
12'd16 : tab = 23'b01111110011101100110000;
12'd17 : tab = 23'b01111110010111101010111;
12'd18 : tab = 23'b01111110010001101111110;
12'd19 : tab = 23'b01111110001011110101001;
12'd20 : tab = 23'b01111110000101111010110;
12'd21 : tab = 23'b01111110000000000000101;
12'd22 : tab = 23'b01111101111010000110101;
12'd23 : tab = 23'b01111101110100001101000;
12'd24 : tab = 23'b01111101101110010011101;
12'd25 : tab = 23'b01111101101000011010100;
12'd26 : tab = 23'b01111101100010100001111;
12'd27 : tab = 23'b01111101011100101001010;
12'd28 : tab = 23'b01111101010110110001000;
12'd29 : tab = 23'b01111101010000111001000;
12'd30 : tab = 23'b01111101001011000001010;
12'd31 : tab = 23'b01111101000101001001110;
12'd32 : tab = 23'b01111100111111010010110;
12'd33 : tab = 23'b01111100111001011011110;
12'd34 : tab = 23'b01111100110011100101010;
12'd35 : tab = 23'b01111100101101101110111;
12'd36 : tab = 23'b01111100100111111000110;
12'd37 : tab = 23'b01111100100010000010110;
12'd38 : tab = 23'b01111100011100001101010;
12'd39 : tab = 23'b01111100010110011000001;
12'd40 : tab = 23'b01111100010000100011000;
12'd41 : tab = 23'b01111100001010101110010;
12'd42 : tab = 23'b01111100000100111001110;
12'd43 : tab = 23'b01111011111111000101100;
12'd44 : tab = 23'b01111011111001010001100;
12'd45 : tab = 23'b01111011110011011110000;
12'd46 : tab = 23'b01111011101101101010011;
12'd47 : tab = 23'b01111011100111110111011;
12'd48 : tab = 23'b01111011100010000100100;
12'd49 : tab = 23'b01111011011100010001111;
12'd50 : tab = 23'b01111011010110011111100;
12'd51 : tab = 23'b01111011010000101101100;
12'd52 : tab = 23'b01111011001010111011110;
12'd53 : tab = 23'b01111011000101001010000;
12'd54 : tab = 23'b01111010111111011000110;
12'd55 : tab = 23'b01111010111001100111101;
12'd56 : tab = 23'b01111010110011110111000;
12'd57 : tab = 23'b01111010101110000110011;
12'd58 : tab = 23'b01111010101000010110000;
12'd59 : tab = 23'b01111010100010100110010;
12'd60 : tab = 23'b01111010011100110110011;
12'd61 : tab = 23'b01111010010111000111000;
12'd62 : tab = 23'b01111010010001010111111;
12'd63 : tab = 23'b01111010001011101000111;
12'd64 : tab = 23'b01111010000101111010010;
12'd65 : tab = 23'b01111010000000001011110;
12'd66 : tab = 23'b01111001111010011101101;
12'd67 : tab = 23'b01111001110100101111110;
12'd68 : tab = 23'b01111001101111000010000;
12'd69 : tab = 23'b01111001101001010100110;
12'd70 : tab = 23'b01111001100011100111101;
12'd71 : tab = 23'b01111001011101111010110;
12'd72 : tab = 23'b01111001011000001110001;
12'd73 : tab = 23'b01111001010010100001110;
12'd74 : tab = 23'b01111001001100110101110;
12'd75 : tab = 23'b01111001000111001001110;
12'd76 : tab = 23'b01111001000001011110011;
12'd77 : tab = 23'b01111000111011110010111;
12'd78 : tab = 23'b01111000110110000111110;
12'd79 : tab = 23'b01111000110000011101001;
12'd80 : tab = 23'b01111000101010110010100;
12'd81 : tab = 23'b01111000100101001000010;
12'd82 : tab = 23'b01111000011111011110010;
12'd83 : tab = 23'b01111000011001110100011;
12'd84 : tab = 23'b01111000010100001010111;
12'd85 : tab = 23'b01111000001110100001100;
12'd86 : tab = 23'b01111000001000111000101;
12'd87 : tab = 23'b01111000000011001111110;
12'd88 : tab = 23'b01110111111101100111010;
12'd89 : tab = 23'b01110111110111111111000;
12'd90 : tab = 23'b01110111110010010111000;
12'd91 : tab = 23'b01110111101100101111001;
12'd92 : tab = 23'b01110111100111000111110;
12'd93 : tab = 23'b01110111100001100000100;
12'd94 : tab = 23'b01110111011011111001100;
12'd95 : tab = 23'b01110111010110010010110;
12'd96 : tab = 23'b01110111010000101100010;
12'd97 : tab = 23'b01110111001011000110000;
12'd98 : tab = 23'b01110111000101100000000;
12'd99 : tab = 23'b01110110111111111010010;
12'd100 : tab = 23'b01110110111010010100110;
12'd101 : tab = 23'b01110110110100101111100;
12'd102 : tab = 23'b01110110101111001010100;
12'd103 : tab = 23'b01110110101001100101110;
12'd104 : tab = 23'b01110110100100000001010;
12'd105 : tab = 23'b01110110011110011101000;
12'd106 : tab = 23'b01110110011000111001000;
12'd107 : tab = 23'b01110110010011010101010;
12'd108 : tab = 23'b01110110001101110001110;
12'd109 : tab = 23'b01110110001000001110100;
12'd110 : tab = 23'b01110110000010101011011;
12'd111 : tab = 23'b01110101111101001000110;
12'd112 : tab = 23'b01110101110111100110001;
12'd113 : tab = 23'b01110101110010000011110;
12'd114 : tab = 23'b01110101101100100001110;
12'd115 : tab = 23'b01110101100111000000000;
12'd116 : tab = 23'b01110101100001011110100;
12'd117 : tab = 23'b01110101011011111101010;
12'd118 : tab = 23'b01110101010110011100001;
12'd119 : tab = 23'b01110101010000111011010;
12'd120 : tab = 23'b01110101001011011010101;
12'd121 : tab = 23'b01110101000101111010100;
12'd122 : tab = 23'b01110101000000011010011;
12'd123 : tab = 23'b01110100111010111010100;
12'd124 : tab = 23'b01110100110101011011000;
12'd125 : tab = 23'b01110100101111111011100;
12'd126 : tab = 23'b01110100101010011100100;
12'd127 : tab = 23'b01110100100100111101110;
12'd128 : tab = 23'b01110100011111011111000;
12'd129 : tab = 23'b01110100011010000000101;
12'd130 : tab = 23'b01110100010100100010100;
12'd131 : tab = 23'b01110100001111000100101;
12'd132 : tab = 23'b01110100001001100111000;
12'd133 : tab = 23'b01110100000100001001100;
12'd134 : tab = 23'b01110011111110101100011;
12'd135 : tab = 23'b01110011111001001111100;
12'd136 : tab = 23'b01110011110011110010110;
12'd137 : tab = 23'b01110011101110010110010;
12'd138 : tab = 23'b01110011101000111010000;
12'd139 : tab = 23'b01110011100011011110001;
12'd140 : tab = 23'b01110011011110000010010;
12'd141 : tab = 23'b01110011011000100110110;
12'd142 : tab = 23'b01110011010011001011100;
12'd143 : tab = 23'b01110011001101110000100;
12'd144 : tab = 23'b01110011001000010101110;
12'd145 : tab = 23'b01110011000010111011010;
12'd146 : tab = 23'b01110010111101100000111;
12'd147 : tab = 23'b01110010111000000110111;
12'd148 : tab = 23'b01110010110010101101000;
12'd149 : tab = 23'b01110010101101010011010;
12'd150 : tab = 23'b01110010100111111010000;
12'd151 : tab = 23'b01110010100010100000111;
12'd152 : tab = 23'b01110010011101001000000;
12'd153 : tab = 23'b01110010010111101111010;
12'd154 : tab = 23'b01110010010010010110110;
12'd155 : tab = 23'b01110010001100111110100;
12'd156 : tab = 23'b01110010000111100110110;
12'd157 : tab = 23'b01110010000010001111000;
12'd158 : tab = 23'b01110001111100110111100;
12'd159 : tab = 23'b01110001110111100000010;
12'd160 : tab = 23'b01110001110010001001010;
12'd161 : tab = 23'b01110001101100110010010;
12'd162 : tab = 23'b01110001100111011011111;
12'd163 : tab = 23'b01110001100010000101100;
12'd164 : tab = 23'b01110001011100101111100;
12'd165 : tab = 23'b01110001010111011001100;
12'd166 : tab = 23'b01110001010010000011111;
12'd167 : tab = 23'b01110001001100101110100;
12'd168 : tab = 23'b01110001000111011001010;
12'd169 : tab = 23'b01110001000010000100011;
12'd170 : tab = 23'b01110000111100101111110;
12'd171 : tab = 23'b01110000110111011011010;
12'd172 : tab = 23'b01110000110010000110111;
12'd173 : tab = 23'b01110000101100110011000;
12'd174 : tab = 23'b01110000100111011111010;
12'd175 : tab = 23'b01110000100010001011101;
12'd176 : tab = 23'b01110000011100111000010;
12'd177 : tab = 23'b01110000010111100101001;
12'd178 : tab = 23'b01110000010010010010010;
12'd179 : tab = 23'b01110000001100111111101;
12'd180 : tab = 23'b01110000000111101101010;
12'd181 : tab = 23'b01110000000010011011000;
12'd182 : tab = 23'b01101111111101001001000;
12'd183 : tab = 23'b01101111110111110111011;
12'd184 : tab = 23'b01101111110010100101111;
12'd185 : tab = 23'b01101111101101010100100;
12'd186 : tab = 23'b01101111101000000011100;
12'd187 : tab = 23'b01101111100010110010110;
12'd188 : tab = 23'b01101111011101100010000;
12'd189 : tab = 23'b01101111011000010001110;
12'd190 : tab = 23'b01101111010011000001100;
12'd191 : tab = 23'b01101111001101110001100;
12'd192 : tab = 23'b01101111001000100010000;
12'd193 : tab = 23'b01101111000011010010100;
12'd194 : tab = 23'b01101110111110000011000;
12'd195 : tab = 23'b01101110111000110100010;
12'd196 : tab = 23'b01101110110011100101010;
12'd197 : tab = 23'b01101110101110010110110;
12'd198 : tab = 23'b01101110101001001000010;
12'd199 : tab = 23'b01101110100011111010010;
12'd200 : tab = 23'b01101110011110101100100;
12'd201 : tab = 23'b01101110011001011110101;
12'd202 : tab = 23'b01101110010100010001010;
12'd203 : tab = 23'b01101110001111000100000;
12'd204 : tab = 23'b01101110001001110111000;
12'd205 : tab = 23'b01101110000100101010000;
12'd206 : tab = 23'b01101101111111011101100;
12'd207 : tab = 23'b01101101111010010001010;
12'd208 : tab = 23'b01101101110101000101000;
12'd209 : tab = 23'b01101101101111111001001;
12'd210 : tab = 23'b01101101101010101101100;
12'd211 : tab = 23'b01101101100101100010000;
12'd212 : tab = 23'b01101101100000010110110;
12'd213 : tab = 23'b01101101011011001011110;
12'd214 : tab = 23'b01101101010110000000110;
12'd215 : tab = 23'b01101101010000110110010;
12'd216 : tab = 23'b01101101001011101011111;
12'd217 : tab = 23'b01101101000110100001101;
12'd218 : tab = 23'b01101101000001010111110;
12'd219 : tab = 23'b01101100111100001110000;
12'd220 : tab = 23'b01101100110111000100100;
12'd221 : tab = 23'b01101100110001111011010;
12'd222 : tab = 23'b01101100101100110010010;
12'd223 : tab = 23'b01101100100111101001011;
12'd224 : tab = 23'b01101100100010100000110;
12'd225 : tab = 23'b01101100011101011000010;
12'd226 : tab = 23'b01101100011000010000000;
12'd227 : tab = 23'b01101100010011001000001;
12'd228 : tab = 23'b01101100001110000000010;
12'd229 : tab = 23'b01101100001000111000110;
12'd230 : tab = 23'b01101100000011110001100;
12'd231 : tab = 23'b01101011111110101010010;
12'd232 : tab = 23'b01101011111001100011100;
12'd233 : tab = 23'b01101011110100011100101;
12'd234 : tab = 23'b01101011101111010110010;
12'd235 : tab = 23'b01101011101010010000000;
12'd236 : tab = 23'b01101011100101001001111;
12'd237 : tab = 23'b01101011100000000100000;
12'd238 : tab = 23'b01101011011010111110100;
12'd239 : tab = 23'b01101011010101111001000;
12'd240 : tab = 23'b01101011010000110011111;
12'd241 : tab = 23'b01101011001011101110111;
12'd242 : tab = 23'b01101011000110101010001;
12'd243 : tab = 23'b01101011000001100101100;
12'd244 : tab = 23'b01101010111100100001010;
12'd245 : tab = 23'b01101010110111011101001;
12'd246 : tab = 23'b01101010110010011001001;
12'd247 : tab = 23'b01101010101101010101100;
12'd248 : tab = 23'b01101010101000010001111;
12'd249 : tab = 23'b01101010100011001110101;
12'd250 : tab = 23'b01101010011110001011110;
12'd251 : tab = 23'b01101010011001001000110;
12'd252 : tab = 23'b01101010010100000110001;
12'd253 : tab = 23'b01101010001111000011101;
12'd254 : tab = 23'b01101010001010000001010;
12'd255 : tab = 23'b01101010000100111111011;
12'd256 : tab = 23'b01101001111111111101101;
12'd257 : tab = 23'b01101001111010111100000;
12'd258 : tab = 23'b01101001110101111010101;
12'd259 : tab = 23'b01101001110000111001011;
12'd260 : tab = 23'b01101001101011111000010;
12'd261 : tab = 23'b01101001100110110111101;
12'd262 : tab = 23'b01101001100001110111000;
12'd263 : tab = 23'b01101001011100110110110;
12'd264 : tab = 23'b01101001010111110110100;
12'd265 : tab = 23'b01101001010010110110110;
12'd266 : tab = 23'b01101001001101110111000;
12'd267 : tab = 23'b01101001001000110111100;
12'd268 : tab = 23'b01101001000011111000001;
12'd269 : tab = 23'b01101000111110111001000;
12'd270 : tab = 23'b01101000111001111010001;
12'd271 : tab = 23'b01101000110100111011011;
12'd272 : tab = 23'b01101000101111111101000;
12'd273 : tab = 23'b01101000101010111110101;
12'd274 : tab = 23'b01101000100110000000101;
12'd275 : tab = 23'b01101000100001000010101;
12'd276 : tab = 23'b01101000011100000101000;
12'd277 : tab = 23'b01101000010111000111100;
12'd278 : tab = 23'b01101000010010001010010;
12'd279 : tab = 23'b01101000001101001101010;
12'd280 : tab = 23'b01101000001000010000011;
12'd281 : tab = 23'b01101000000011010011110;
12'd282 : tab = 23'b01100111111110010111010;
12'd283 : tab = 23'b01100111111001011011000;
12'd284 : tab = 23'b01100111110100011111000;
12'd285 : tab = 23'b01100111101111100011010;
12'd286 : tab = 23'b01100111101010100111101;
12'd287 : tab = 23'b01100111100101101100001;
12'd288 : tab = 23'b01100111100000110001000;
12'd289 : tab = 23'b01100111011011110101111;
12'd290 : tab = 23'b01100111010110111011000;
12'd291 : tab = 23'b01100111010010000000100;
12'd292 : tab = 23'b01100111001101000110000;
12'd293 : tab = 23'b01100111001000001011111;
12'd294 : tab = 23'b01100111000011010001111;
12'd295 : tab = 23'b01100110111110011000000;
12'd296 : tab = 23'b01100110111001011110011;
12'd297 : tab = 23'b01100110110100100101000;
12'd298 : tab = 23'b01100110101111101011110;
12'd299 : tab = 23'b01100110101010110010110;
12'd300 : tab = 23'b01100110100101111010000;
12'd301 : tab = 23'b01100110100001000001011;
12'd302 : tab = 23'b01100110011100001000111;
12'd303 : tab = 23'b01100110010111010000110;
12'd304 : tab = 23'b01100110010010011000110;
12'd305 : tab = 23'b01100110001101100001000;
12'd306 : tab = 23'b01100110001000101001011;
12'd307 : tab = 23'b01100110000011110001111;
12'd308 : tab = 23'b01100101111110111010101;
12'd309 : tab = 23'b01100101111010000011110;
12'd310 : tab = 23'b01100101110101001100110;
12'd311 : tab = 23'b01100101110000010110010;
12'd312 : tab = 23'b01100101101011011111110;
12'd313 : tab = 23'b01100101100110101001101;
12'd314 : tab = 23'b01100101100001110011100;
12'd315 : tab = 23'b01100101011100111101101;
12'd316 : tab = 23'b01100101011000001000000;
12'd317 : tab = 23'b01100101010011010010110;
12'd318 : tab = 23'b01100101001110011101010;
12'd319 : tab = 23'b01100101001001101000010;
12'd320 : tab = 23'b01100101000100110011100;
12'd321 : tab = 23'b01100100111111111110111;
12'd322 : tab = 23'b01100100111011001010100;
12'd323 : tab = 23'b01100100110110010110000;
12'd324 : tab = 23'b01100100110001100010000;
12'd325 : tab = 23'b01100100101100101110000;
12'd326 : tab = 23'b01100100100111111010011;
12'd327 : tab = 23'b01100100100011000111000;
12'd328 : tab = 23'b01100100011110010011100;
12'd329 : tab = 23'b01100100011001100000101;
12'd330 : tab = 23'b01100100010100101101101;
12'd331 : tab = 23'b01100100001111111011000;
12'd332 : tab = 23'b01100100001011001000011;
12'd333 : tab = 23'b01100100000110010110001;
12'd334 : tab = 23'b01100100000001100100000;
12'd335 : tab = 23'b01100011111100110010000;
12'd336 : tab = 23'b01100011111000000000010;
12'd337 : tab = 23'b01100011110011001110110;
12'd338 : tab = 23'b01100011101110011101010;
12'd339 : tab = 23'b01100011101001101100010;
12'd340 : tab = 23'b01100011100100111011010;
12'd341 : tab = 23'b01100011100000001010011;
12'd342 : tab = 23'b01100011011011011001110;
12'd343 : tab = 23'b01100011010110101001010;
12'd344 : tab = 23'b01100011010001111001010;
12'd345 : tab = 23'b01100011001101001001000;
12'd346 : tab = 23'b01100011001000011001010;
12'd347 : tab = 23'b01100011000011101001110;
12'd348 : tab = 23'b01100010111110111010010;
12'd349 : tab = 23'b01100010111010001010111;
12'd350 : tab = 23'b01100010110101011011110;
12'd351 : tab = 23'b01100010110000101101000;
12'd352 : tab = 23'b01100010101011111110010;
12'd353 : tab = 23'b01100010100111001111110;
12'd354 : tab = 23'b01100010100010100001100;
12'd355 : tab = 23'b01100010011101110011100;
12'd356 : tab = 23'b01100010011001000101011;
12'd357 : tab = 23'b01100010010100010111101;
12'd358 : tab = 23'b01100010001111101010000;
12'd359 : tab = 23'b01100010001010111100110;
12'd360 : tab = 23'b01100010000110001111011;
12'd361 : tab = 23'b01100010000001100010100;
12'd362 : tab = 23'b01100001111100110101110;
12'd363 : tab = 23'b01100001111000001001001;
12'd364 : tab = 23'b01100001110011011100100;
12'd365 : tab = 23'b01100001101110110000010;
12'd366 : tab = 23'b01100001101010000100010;
12'd367 : tab = 23'b01100001100101011000011;
12'd368 : tab = 23'b01100001100000101100110;
12'd369 : tab = 23'b01100001011100000001010;
12'd370 : tab = 23'b01100001010111010101111;
12'd371 : tab = 23'b01100001010010101010101;
12'd372 : tab = 23'b01100001001101111111110;
12'd373 : tab = 23'b01100001001001010101000;
12'd374 : tab = 23'b01100001000100101010011;
12'd375 : tab = 23'b01100000111111111111111;
12'd376 : tab = 23'b01100000111011010101110;
12'd377 : tab = 23'b01100000110110101011110;
12'd378 : tab = 23'b01100000110010000010000;
12'd379 : tab = 23'b01100000101101011000010;
12'd380 : tab = 23'b01100000101000101110110;
12'd381 : tab = 23'b01100000100100000101011;
12'd382 : tab = 23'b01100000011111011100011;
12'd383 : tab = 23'b01100000011010110011100;
12'd384 : tab = 23'b01100000010110001010110;
12'd385 : tab = 23'b01100000010001100010001;
12'd386 : tab = 23'b01100000001100111001110;
12'd387 : tab = 23'b01100000001000010001100;
12'd388 : tab = 23'b01100000000011101001100;
12'd389 : tab = 23'b01011111111111000001110;
12'd390 : tab = 23'b01011111111010011010010;
12'd391 : tab = 23'b01011111110101110010101;
12'd392 : tab = 23'b01011111110001001011011;
12'd393 : tab = 23'b01011111101100100100010;
12'd394 : tab = 23'b01011111100111111101010;
12'd395 : tab = 23'b01011111100011010110100;
12'd396 : tab = 23'b01011111011110110000001;
12'd397 : tab = 23'b01011111011010001001101;
12'd398 : tab = 23'b01011111010101100011100;
12'd399 : tab = 23'b01011111010000111101100;
12'd400 : tab = 23'b01011111001100010111101;
12'd401 : tab = 23'b01011111000111110001111;
12'd402 : tab = 23'b01011111000011001100011;
12'd403 : tab = 23'b01011110111110100111001;
12'd404 : tab = 23'b01011110111010000010000;
12'd405 : tab = 23'b01011110110101011101001;
12'd406 : tab = 23'b01011110110000111000010;
12'd407 : tab = 23'b01011110101100010011110;
12'd408 : tab = 23'b01011110100111101111010;
12'd409 : tab = 23'b01011110100011001011000;
12'd410 : tab = 23'b01011110011110100111000;
12'd411 : tab = 23'b01011110011010000011001;
12'd412 : tab = 23'b01011110010101011111011;
12'd413 : tab = 23'b01011110010000111100000;
12'd414 : tab = 23'b01011110001100011000101;
12'd415 : tab = 23'b01011110000111110101100;
12'd416 : tab = 23'b01011110000011010010100;
12'd417 : tab = 23'b01011101111110101111110;
12'd418 : tab = 23'b01011101111010001101000;
12'd419 : tab = 23'b01011101110101101010100;
12'd420 : tab = 23'b01011101110001001000010;
12'd421 : tab = 23'b01011101101100100110010;
12'd422 : tab = 23'b01011101101000000100011;
12'd423 : tab = 23'b01011101100011100010100;
12'd424 : tab = 23'b01011101011111000001000;
12'd425 : tab = 23'b01011101011010011111110;
12'd426 : tab = 23'b01011101010101111110100;
12'd427 : tab = 23'b01011101010001011101010;
12'd428 : tab = 23'b01011101001100111100100;
12'd429 : tab = 23'b01011101001000011011110;
12'd430 : tab = 23'b01011101000011111011010;
12'd431 : tab = 23'b01011100111111011010111;
12'd432 : tab = 23'b01011100111010111010110;
12'd433 : tab = 23'b01011100110110011010110;
12'd434 : tab = 23'b01011100110001111011000;
12'd435 : tab = 23'b01011100101101011011010;
12'd436 : tab = 23'b01011100101000111011111;
12'd437 : tab = 23'b01011100100100011100100;
12'd438 : tab = 23'b01011100011111111101011;
12'd439 : tab = 23'b01011100011011011110100;
12'd440 : tab = 23'b01011100010110111111110;
12'd441 : tab = 23'b01011100010010100001000;
12'd442 : tab = 23'b01011100001110000010101;
12'd443 : tab = 23'b01011100001001100100011;
12'd444 : tab = 23'b01011100000101000110010;
12'd445 : tab = 23'b01011100000000101000010;
12'd446 : tab = 23'b01011011111100001010100;
12'd447 : tab = 23'b01011011110111101101000;
12'd448 : tab = 23'b01011011110011001111101;
12'd449 : tab = 23'b01011011101110110010011;
12'd450 : tab = 23'b01011011101010010101010;
12'd451 : tab = 23'b01011011100101111000100;
12'd452 : tab = 23'b01011011100001011011110;
12'd453 : tab = 23'b01011011011100111111010;
12'd454 : tab = 23'b01011011011000100010110;
12'd455 : tab = 23'b01011011010100000110101;
12'd456 : tab = 23'b01011011001111101010100;
12'd457 : tab = 23'b01011011001011001110101;
12'd458 : tab = 23'b01011011000110110011000;
12'd459 : tab = 23'b01011011000010010111100;
12'd460 : tab = 23'b01011010111101111100000;
12'd461 : tab = 23'b01011010111001100001000;
12'd462 : tab = 23'b01011010110101000101110;
12'd463 : tab = 23'b01011010110000101011000;
12'd464 : tab = 23'b01011010101100010000010;
12'd465 : tab = 23'b01011010100111110101111;
12'd466 : tab = 23'b01011010100011011011011;
12'd467 : tab = 23'b01011010011111000001011;
12'd468 : tab = 23'b01011010011010100111010;
12'd469 : tab = 23'b01011010010110001101100;
12'd470 : tab = 23'b01011010010001110011110;
12'd471 : tab = 23'b01011010001101011010010;
12'd472 : tab = 23'b01011010001001000000111;
12'd473 : tab = 23'b01011010000100100111110;
12'd474 : tab = 23'b01011010000000001110110;
12'd475 : tab = 23'b01011001111011110101111;
12'd476 : tab = 23'b01011001110111011101010;
12'd477 : tab = 23'b01011001110011000100111;
12'd478 : tab = 23'b01011001101110101100100;
12'd479 : tab = 23'b01011001101010010100010;
12'd480 : tab = 23'b01011001100101111100010;
12'd481 : tab = 23'b01011001100001100100011;
12'd482 : tab = 23'b01011001011101001100110;
12'd483 : tab = 23'b01011001011000110101010;
12'd484 : tab = 23'b01011001010100011101111;
12'd485 : tab = 23'b01011001010000000110110;
12'd486 : tab = 23'b01011001001011101111110;
12'd487 : tab = 23'b01011001000111011000111;
12'd488 : tab = 23'b01011001000011000010010;
12'd489 : tab = 23'b01011000111110101011110;
12'd490 : tab = 23'b01011000111010010101011;
12'd491 : tab = 23'b01011000110101111111010;
12'd492 : tab = 23'b01011000110001101001010;
12'd493 : tab = 23'b01011000101101010011011;
12'd494 : tab = 23'b01011000101000111101101;
12'd495 : tab = 23'b01011000100100101000000;
12'd496 : tab = 23'b01011000100000010010110;
12'd497 : tab = 23'b01011000011011111101100;
12'd498 : tab = 23'b01011000010111101000100;
12'd499 : tab = 23'b01011000010011010011110;
12'd500 : tab = 23'b01011000001110111111000;
12'd501 : tab = 23'b01011000001010101010010;
12'd502 : tab = 23'b01011000000110010110000;
12'd503 : tab = 23'b01011000000010000001110;
12'd504 : tab = 23'b01010111111101101101101;
12'd505 : tab = 23'b01010111111001011001110;
12'd506 : tab = 23'b01010111110101000110000;
12'd507 : tab = 23'b01010111110000110010100;
12'd508 : tab = 23'b01010111101100011111001;
12'd509 : tab = 23'b01010111101000001011110;
12'd510 : tab = 23'b01010111100011111000110;
12'd511 : tab = 23'b01010111011111100101111;
12'd512 : tab = 23'b01010111011011010011000;
12'd513 : tab = 23'b01010111010111000000100;
12'd514 : tab = 23'b01010111010010101101111;
12'd515 : tab = 23'b01010111001110011011101;
12'd516 : tab = 23'b01010111001010001001101;
12'd517 : tab = 23'b01010111000101110111101;
12'd518 : tab = 23'b01010111000001100101110;
12'd519 : tab = 23'b01010110111101010100010;
12'd520 : tab = 23'b01010110111001000010101;
12'd521 : tab = 23'b01010110110100110001100;
12'd522 : tab = 23'b01010110110000100000010;
12'd523 : tab = 23'b01010110101100001111001;
12'd524 : tab = 23'b01010110100111111110010;
12'd525 : tab = 23'b01010110100011101101101;
12'd526 : tab = 23'b01010110011111011101001;
12'd527 : tab = 23'b01010110011011001100110;
12'd528 : tab = 23'b01010110010110111100100;
12'd529 : tab = 23'b01010110010010101100100;
12'd530 : tab = 23'b01010110001110011100100;
12'd531 : tab = 23'b01010110001010001100111;
12'd532 : tab = 23'b01010110000101111101011;
12'd533 : tab = 23'b01010110000001101101110;
12'd534 : tab = 23'b01010101111101011110100;
12'd535 : tab = 23'b01010101111001001111100;
12'd536 : tab = 23'b01010101110101000000100;
12'd537 : tab = 23'b01010101110000110001101;
12'd538 : tab = 23'b01010101101100100011000;
12'd539 : tab = 23'b01010101101000010100101;
12'd540 : tab = 23'b01010101100100000110010;
12'd541 : tab = 23'b01010101011111111000000;
12'd542 : tab = 23'b01010101011011101010000;
12'd543 : tab = 23'b01010101010111011100010;
12'd544 : tab = 23'b01010101010011001110100;
12'd545 : tab = 23'b01010101001111000001000;
12'd546 : tab = 23'b01010101001010110011101;
12'd547 : tab = 23'b01010101000110100110010;
12'd548 : tab = 23'b01010101000010011001011;
12'd549 : tab = 23'b01010100111110001100011;
12'd550 : tab = 23'b01010100111001111111110;
12'd551 : tab = 23'b01010100110101110011000;
12'd552 : tab = 23'b01010100110001100110110;
12'd553 : tab = 23'b01010100101101011010011;
12'd554 : tab = 23'b01010100101001001110001;
12'd555 : tab = 23'b01010100100101000010001;
12'd556 : tab = 23'b01010100100000110110010;
12'd557 : tab = 23'b01010100011100101010101;
12'd558 : tab = 23'b01010100011000011111000;
12'd559 : tab = 23'b01010100010100010011110;
12'd560 : tab = 23'b01010100010000001000100;
12'd561 : tab = 23'b01010100001011111101100;
12'd562 : tab = 23'b01010100000111110010101;
12'd563 : tab = 23'b01010100000011100111111;
12'd564 : tab = 23'b01010011111111011101010;
12'd565 : tab = 23'b01010011111011010010110;
12'd566 : tab = 23'b01010011110111001000100;
12'd567 : tab = 23'b01010011110010111110010;
12'd568 : tab = 23'b01010011101110110100100;
12'd569 : tab = 23'b01010011101010101010100;
12'd570 : tab = 23'b01010011100110100000111;
12'd571 : tab = 23'b01010011100010010111010;
12'd572 : tab = 23'b01010011011110001101111;
12'd573 : tab = 23'b01010011011010000100101;
12'd574 : tab = 23'b01010011010101111011101;
12'd575 : tab = 23'b01010011010001110010110;
12'd576 : tab = 23'b01010011001101101001111;
12'd577 : tab = 23'b01010011001001100001010;
12'd578 : tab = 23'b01010011000101011000110;
12'd579 : tab = 23'b01010011000001010000100;
12'd580 : tab = 23'b01010010111101001000010;
12'd581 : tab = 23'b01010010111001000000010;
12'd582 : tab = 23'b01010010110100111000011;
12'd583 : tab = 23'b01010010110000110000101;
12'd584 : tab = 23'b01010010101100101001001;
12'd585 : tab = 23'b01010010101000100001110;
12'd586 : tab = 23'b01010010100100011010011;
12'd587 : tab = 23'b01010010100000010011010;
12'd588 : tab = 23'b01010010011100001100011;
12'd589 : tab = 23'b01010010011000000101100;
12'd590 : tab = 23'b01010010010011111110110;
12'd591 : tab = 23'b01010010001111111000010;
12'd592 : tab = 23'b01010010001011110001111;
12'd593 : tab = 23'b01010010000111101011110;
12'd594 : tab = 23'b01010010000011100101100;
12'd595 : tab = 23'b01010001111111011111101;
12'd596 : tab = 23'b01010001111011011001111;
12'd597 : tab = 23'b01010001110111010100010;
12'd598 : tab = 23'b01010001110011001110111;
12'd599 : tab = 23'b01010001101111001001011;
12'd600 : tab = 23'b01010001101011000100010;
12'd601 : tab = 23'b01010001100110111111010;
12'd602 : tab = 23'b01010001100010111010011;
12'd603 : tab = 23'b01010001011110110101100;
12'd604 : tab = 23'b01010001011010110001000;
12'd605 : tab = 23'b01010001010110101100100;
12'd606 : tab = 23'b01010001010010101000010;
12'd607 : tab = 23'b01010001001110100100001;
12'd608 : tab = 23'b01010001001010100000001;
12'd609 : tab = 23'b01010001000110011100010;
12'd610 : tab = 23'b01010001000010011000100;
12'd611 : tab = 23'b01010000111110010101000;
12'd612 : tab = 23'b01010000111010010001100;
12'd613 : tab = 23'b01010000110110001110010;
12'd614 : tab = 23'b01010000110010001011001;
12'd615 : tab = 23'b01010000101110001000010;
12'd616 : tab = 23'b01010000101010000101011;
12'd617 : tab = 23'b01010000100110000010110;
12'd618 : tab = 23'b01010000100010000000001;
12'd619 : tab = 23'b01010000011101111101100;
12'd620 : tab = 23'b01010000011001111011011;
12'd621 : tab = 23'b01010000010101111001011;
12'd622 : tab = 23'b01010000010001110111011;
12'd623 : tab = 23'b01010000001101110101100;
12'd624 : tab = 23'b01010000001001110011111;
12'd625 : tab = 23'b01010000000101110010010;
12'd626 : tab = 23'b01010000000001110000111;
12'd627 : tab = 23'b01001111111101101111101;
12'd628 : tab = 23'b01001111111001101110100;
12'd629 : tab = 23'b01001111110101101101110;
12'd630 : tab = 23'b01001111110001101100110;
12'd631 : tab = 23'b01001111101101101100001;
12'd632 : tab = 23'b01001111101001101011101;
12'd633 : tab = 23'b01001111100101101011010;
12'd634 : tab = 23'b01001111100001101011000;
12'd635 : tab = 23'b01001111011101101011000;
12'd636 : tab = 23'b01001111011001101011000;
12'd637 : tab = 23'b01001111010101101011010;
12'd638 : tab = 23'b01001111010001101011100;
12'd639 : tab = 23'b01001111001101101100000;
12'd640 : tab = 23'b01001111001001101100101;
12'd641 : tab = 23'b01001111000101101101011;
12'd642 : tab = 23'b01001111000001101110010;
12'd643 : tab = 23'b01001110111101101111011;
12'd644 : tab = 23'b01001110111001110000100;
12'd645 : tab = 23'b01001110110101110001111;
12'd646 : tab = 23'b01001110110001110011010;
12'd647 : tab = 23'b01001110101101110101000;
12'd648 : tab = 23'b01001110101001110110110;
12'd649 : tab = 23'b01001110100101111000110;
12'd650 : tab = 23'b01001110100001111010101;
12'd651 : tab = 23'b01001110011101111100111;
12'd652 : tab = 23'b01001110011001111111000;
12'd653 : tab = 23'b01001110010110000001100;
12'd654 : tab = 23'b01001110010010000100010;
12'd655 : tab = 23'b01001110001110000111000;
12'd656 : tab = 23'b01001110001010001001110;
12'd657 : tab = 23'b01001110000110001100111;
12'd658 : tab = 23'b01001110000010010000000;
12'd659 : tab = 23'b01001101111110010011011;
12'd660 : tab = 23'b01001101111010010110110;
12'd661 : tab = 23'b01001101110110011010100;
12'd662 : tab = 23'b01001101110010011110000;
12'd663 : tab = 23'b01001101101110100010000;
12'd664 : tab = 23'b01001101101010100110000;
12'd665 : tab = 23'b01001101100110101010010;
12'd666 : tab = 23'b01001101100010101110100;
12'd667 : tab = 23'b01001101011110110010110;
12'd668 : tab = 23'b01001101011010110111011;
12'd669 : tab = 23'b01001101010110111100001;
12'd670 : tab = 23'b01001101010011000001000;
12'd671 : tab = 23'b01001101001111000101111;
12'd672 : tab = 23'b01001101001011001011000;
12'd673 : tab = 23'b01001101000111010000010;
12'd674 : tab = 23'b01001101000011010101110;
12'd675 : tab = 23'b01001100111111011011010;
12'd676 : tab = 23'b01001100111011100001000;
12'd677 : tab = 23'b01001100110111100110110;
12'd678 : tab = 23'b01001100110011101100110;
12'd679 : tab = 23'b01001100101111110010110;
12'd680 : tab = 23'b01001100101011111001000;
12'd681 : tab = 23'b01001100100111111111010;
12'd682 : tab = 23'b01001100100100000101110;
12'd683 : tab = 23'b01001100100000001100100;
12'd684 : tab = 23'b01001100011100010011010;
12'd685 : tab = 23'b01001100011000011010001;
12'd686 : tab = 23'b01001100010100100001010;
12'd687 : tab = 23'b01001100010000101000010;
12'd688 : tab = 23'b01001100001100101111110;
12'd689 : tab = 23'b01001100001000110111000;
12'd690 : tab = 23'b01001100000100111110101;
12'd691 : tab = 23'b01001100000001000110011;
12'd692 : tab = 23'b01001011111101001110010;
12'd693 : tab = 23'b01001011111001010110010;
12'd694 : tab = 23'b01001011110101011110011;
12'd695 : tab = 23'b01001011110001100110110;
12'd696 : tab = 23'b01001011101101101111000;
12'd697 : tab = 23'b01001011101001110111101;
12'd698 : tab = 23'b01001011100110000000010;
12'd699 : tab = 23'b01001011100010001001000;
12'd700 : tab = 23'b01001011011110010010000;
12'd701 : tab = 23'b01001011011010011011001;
12'd702 : tab = 23'b01001011010110100100010;
12'd703 : tab = 23'b01001011010010101101110;
12'd704 : tab = 23'b01001011001110110111001;
12'd705 : tab = 23'b01001011001011000000110;
12'd706 : tab = 23'b01001011000111001010011;
12'd707 : tab = 23'b01001011000011010100010;
12'd708 : tab = 23'b01001010111111011110011;
12'd709 : tab = 23'b01001010111011101000100;
12'd710 : tab = 23'b01001010110111110010110;
12'd711 : tab = 23'b01001010110011111101010;
12'd712 : tab = 23'b01001010110000000111110;
12'd713 : tab = 23'b01001010101100010010100;
12'd714 : tab = 23'b01001010101000011101010;
12'd715 : tab = 23'b01001010100100101000010;
12'd716 : tab = 23'b01001010100000110011010;
12'd717 : tab = 23'b01001010011100111110100;
12'd718 : tab = 23'b01001010011001001001111;
12'd719 : tab = 23'b01001010010101010101011;
12'd720 : tab = 23'b01001010010001100000111;
12'd721 : tab = 23'b01001010001101101100101;
12'd722 : tab = 23'b01001010001001111000100;
12'd723 : tab = 23'b01001010000110000100100;
12'd724 : tab = 23'b01001010000010010000110;
12'd725 : tab = 23'b01001001111110011101000;
12'd726 : tab = 23'b01001001111010101001011;
12'd727 : tab = 23'b01001001110110110110000;
12'd728 : tab = 23'b01001001110011000010110;
12'd729 : tab = 23'b01001001101111001111100;
12'd730 : tab = 23'b01001001101011011100010;
12'd731 : tab = 23'b01001001100111101001011;
12'd732 : tab = 23'b01001001100011110110110;
12'd733 : tab = 23'b01001001100000000011111;
12'd734 : tab = 23'b01001001011100010001011;
12'd735 : tab = 23'b01001001011000011111000;
12'd736 : tab = 23'b01001001010100101100110;
12'd737 : tab = 23'b01001001010000111010100;
12'd738 : tab = 23'b01001001001101001000100;
12'd739 : tab = 23'b01001001001001010110100;
12'd740 : tab = 23'b01001001000101100100111;
12'd741 : tab = 23'b01001001000001110011010;
12'd742 : tab = 23'b01001000111110000001110;
12'd743 : tab = 23'b01001000111010010000011;
12'd744 : tab = 23'b01001000110110011111000;
12'd745 : tab = 23'b01001000110010101110000;
12'd746 : tab = 23'b01001000101110111101000;
12'd747 : tab = 23'b01001000101011001100010;
12'd748 : tab = 23'b01001000100111011011011;
12'd749 : tab = 23'b01001000100011101011000;
12'd750 : tab = 23'b01001000011111111010011;
12'd751 : tab = 23'b01001000011100001010000;
12'd752 : tab = 23'b01001000011000011001110;
12'd753 : tab = 23'b01001000010100101001110;
12'd754 : tab = 23'b01001000010000111001110;
12'd755 : tab = 23'b01001000001101001001111;
12'd756 : tab = 23'b01001000001001011010010;
12'd757 : tab = 23'b01001000000101101010110;
12'd758 : tab = 23'b01001000000001111011010;
12'd759 : tab = 23'b01000111111110001100000;
12'd760 : tab = 23'b01000111111010011100110;
12'd761 : tab = 23'b01000111110110101101110;
12'd762 : tab = 23'b01000111110010111110110;
12'd763 : tab = 23'b01000111101111010000000;
12'd764 : tab = 23'b01000111101011100001010;
12'd765 : tab = 23'b01000111100111110010110;
12'd766 : tab = 23'b01000111100100000100010;
12'd767 : tab = 23'b01000111100000010110001;
12'd768 : tab = 23'b01000111011100100111111;
12'd769 : tab = 23'b01000111011000111001111;
12'd770 : tab = 23'b01000111010101001100000;
12'd771 : tab = 23'b01000111010001011110010;
12'd772 : tab = 23'b01000111001101110000101;
12'd773 : tab = 23'b01000111001010000011000;
12'd774 : tab = 23'b01000111000110010101100;
12'd775 : tab = 23'b01000111000010101000010;
12'd776 : tab = 23'b01000110111110111011010;
12'd777 : tab = 23'b01000110111011001110010;
12'd778 : tab = 23'b01000110110111100001010;
12'd779 : tab = 23'b01000110110011110100011;
12'd780 : tab = 23'b01000110110000000111110;
12'd781 : tab = 23'b01000110101100011011010;
12'd782 : tab = 23'b01000110101000101110111;
12'd783 : tab = 23'b01000110100101000010101;
12'd784 : tab = 23'b01000110100001010110011;
12'd785 : tab = 23'b01000110011101101010100;
12'd786 : tab = 23'b01000110011001111110100;
12'd787 : tab = 23'b01000110010110010010110;
12'd788 : tab = 23'b01000110010010100111000;
12'd789 : tab = 23'b01000110001110111011100;
12'd790 : tab = 23'b01000110001011010000001;
12'd791 : tab = 23'b01000110000111100101000;
12'd792 : tab = 23'b01000110000011111001110;
12'd793 : tab = 23'b01000110000000001110110;
12'd794 : tab = 23'b01000101111100100011110;
12'd795 : tab = 23'b01000101111000111001000;
12'd796 : tab = 23'b01000101110101001110100;
12'd797 : tab = 23'b01000101110001100011110;
12'd798 : tab = 23'b01000101101101111001100;
12'd799 : tab = 23'b01000101101010001111001;
12'd800 : tab = 23'b01000101100110100101000;
12'd801 : tab = 23'b01000101100010111011000;
12'd802 : tab = 23'b01000101011111010001000;
12'd803 : tab = 23'b01000101011011100111010;
12'd804 : tab = 23'b01000101010111111101101;
12'd805 : tab = 23'b01000101010100010100000;
12'd806 : tab = 23'b01000101010000101010101;
12'd807 : tab = 23'b01000101001101000001010;
12'd808 : tab = 23'b01000101001001011000001;
12'd809 : tab = 23'b01000101000101101111000;
12'd810 : tab = 23'b01000101000010000110010;
12'd811 : tab = 23'b01000100111110011101010;
12'd812 : tab = 23'b01000100111010110100101;
12'd813 : tab = 23'b01000100110111001100000;
12'd814 : tab = 23'b01000100110011100011101;
12'd815 : tab = 23'b01000100101111111011010;
12'd816 : tab = 23'b01000100101100010011001;
12'd817 : tab = 23'b01000100101000101011000;
12'd818 : tab = 23'b01000100100101000011000;
12'd819 : tab = 23'b01000100100001011011010;
12'd820 : tab = 23'b01000100011101110011100;
12'd821 : tab = 23'b01000100011010001011111;
12'd822 : tab = 23'b01000100010110100100011;
12'd823 : tab = 23'b01000100010010111101001;
12'd824 : tab = 23'b01000100001111010101111;
12'd825 : tab = 23'b01000100001011101110110;
12'd826 : tab = 23'b01000100001000000111110;
12'd827 : tab = 23'b01000100000100100000111;
12'd828 : tab = 23'b01000100000000111010001;
12'd829 : tab = 23'b01000011111101010011100;
12'd830 : tab = 23'b01000011111001101100111;
12'd831 : tab = 23'b01000011110110000110101;
12'd832 : tab = 23'b01000011110010100000011;
12'd833 : tab = 23'b01000011101110111010010;
12'd834 : tab = 23'b01000011101011010100000;
12'd835 : tab = 23'b01000011100111101110010;
12'd836 : tab = 23'b01000011100100001000100;
12'd837 : tab = 23'b01000011100000100010110;
12'd838 : tab = 23'b01000011011100111101010;
12'd839 : tab = 23'b01000011011001010111110;
12'd840 : tab = 23'b01000011010101110010100;
12'd841 : tab = 23'b01000011010010001101010;
12'd842 : tab = 23'b01000011001110101000001;
12'd843 : tab = 23'b01000011001011000011001;
12'd844 : tab = 23'b01000011000111011110011;
12'd845 : tab = 23'b01000011000011111001101;
12'd846 : tab = 23'b01000011000000010101000;
12'd847 : tab = 23'b01000010111100110000101;
12'd848 : tab = 23'b01000010111001001100010;
12'd849 : tab = 23'b01000010110101101000000;
12'd850 : tab = 23'b01000010110010000100000;
12'd851 : tab = 23'b01000010101110011111110;
12'd852 : tab = 23'b01000010101010111100000;
12'd853 : tab = 23'b01000010100111011000010;
12'd854 : tab = 23'b01000010100011110100100;
12'd855 : tab = 23'b01000010100000010001000;
12'd856 : tab = 23'b01000010011100101101101;
12'd857 : tab = 23'b01000010011001001010010;
12'd858 : tab = 23'b01000010010101100111001;
12'd859 : tab = 23'b01000010010010000100000;
12'd860 : tab = 23'b01000010001110100001000;
12'd861 : tab = 23'b01000010001010111110010;
12'd862 : tab = 23'b01000010000111011011100;
12'd863 : tab = 23'b01000010000011111001000;
12'd864 : tab = 23'b01000010000000010110100;
12'd865 : tab = 23'b01000001111100110100000;
12'd866 : tab = 23'b01000001111001010001110;
12'd867 : tab = 23'b01000001110101101111110;
12'd868 : tab = 23'b01000001110010001101101;
12'd869 : tab = 23'b01000001101110101011110;
12'd870 : tab = 23'b01000001101011001010000;
12'd871 : tab = 23'b01000001100111101000010;
12'd872 : tab = 23'b01000001100100000110110;
12'd873 : tab = 23'b01000001100000100101011;
12'd874 : tab = 23'b01000001011101000011111;
12'd875 : tab = 23'b01000001011001100010110;
12'd876 : tab = 23'b01000001010110000001101;
12'd877 : tab = 23'b01000001010010100000110;
12'd878 : tab = 23'b01000001001110111111110;
12'd879 : tab = 23'b01000001001011011111000;
12'd880 : tab = 23'b01000001000111111110100;
12'd881 : tab = 23'b01000001000100011101111;
12'd882 : tab = 23'b01000001000000111101100;
12'd883 : tab = 23'b01000000111101011101010;
12'd884 : tab = 23'b01000000111001111101001;
12'd885 : tab = 23'b01000000110110011101001;
12'd886 : tab = 23'b01000000110010111101000;
12'd887 : tab = 23'b01000000101111011101010;
12'd888 : tab = 23'b01000000101011111101100;
12'd889 : tab = 23'b01000000101000011101110;
12'd890 : tab = 23'b01000000100100111110011;
12'd891 : tab = 23'b01000000100001011111001;
12'd892 : tab = 23'b01000000011101111111111;
12'd893 : tab = 23'b01000000011010100000101;
12'd894 : tab = 23'b01000000010111000001101;
12'd895 : tab = 23'b01000000010011100010110;
12'd896 : tab = 23'b01000000010000000100000;
12'd897 : tab = 23'b01000000001100100101010;
12'd898 : tab = 23'b01000000001001000110101;
12'd899 : tab = 23'b01000000000101101000001;
12'd900 : tab = 23'b01000000000010001001111;
12'd901 : tab = 23'b00111111111110101011101;
12'd902 : tab = 23'b00111111111011001101100;
12'd903 : tab = 23'b00111111110111101111100;
12'd904 : tab = 23'b00111111110100010001100;
12'd905 : tab = 23'b00111111110000110011111;
12'd906 : tab = 23'b00111111101101010110000;
12'd907 : tab = 23'b00111111101001111000101;
12'd908 : tab = 23'b00111111100110011011000;
12'd909 : tab = 23'b00111111100010111101110;
12'd910 : tab = 23'b00111111011111100000100;
12'd911 : tab = 23'b00111111011100000011100;
12'd912 : tab = 23'b00111111011000100110100;
12'd913 : tab = 23'b00111111010101001001101;
12'd914 : tab = 23'b00111111010001101100110;
12'd915 : tab = 23'b00111111001110010000001;
12'd916 : tab = 23'b00111111001010110011100;
12'd917 : tab = 23'b00111111000111010111001;
12'd918 : tab = 23'b00111111000011111010110;
12'd919 : tab = 23'b00111111000000011110100;
12'd920 : tab = 23'b00111110111101000010100;
12'd921 : tab = 23'b00111110111001100110100;
12'd922 : tab = 23'b00111110110110001010101;
12'd923 : tab = 23'b00111110110010101111000;
12'd924 : tab = 23'b00111110101111010011010;
12'd925 : tab = 23'b00111110101011110111101;
12'd926 : tab = 23'b00111110101000011100010;
12'd927 : tab = 23'b00111110100101000000111;
12'd928 : tab = 23'b00111110100001100101110;
12'd929 : tab = 23'b00111110011110001010100;
12'd930 : tab = 23'b00111110011010101111100;
12'd931 : tab = 23'b00111110010111010100110;
12'd932 : tab = 23'b00111110010011111001111;
12'd933 : tab = 23'b00111110010000011111010;
12'd934 : tab = 23'b00111110001101000100101;
12'd935 : tab = 23'b00111110001001101010010;
12'd936 : tab = 23'b00111110000110010000000;
12'd937 : tab = 23'b00111110000010110101110;
12'd938 : tab = 23'b00111101111111011011100;
12'd939 : tab = 23'b00111101111100000001100;
12'd940 : tab = 23'b00111101111000100111100;
12'd941 : tab = 23'b00111101110101001101110;
12'd942 : tab = 23'b00111101110001110100001;
12'd943 : tab = 23'b00111101101110011010100;
12'd944 : tab = 23'b00111101101011000001001;
12'd945 : tab = 23'b00111101100111100111110;
12'd946 : tab = 23'b00111101100100001110100;
12'd947 : tab = 23'b00111101100000110101011;
12'd948 : tab = 23'b00111101011101011100011;
12'd949 : tab = 23'b00111101011010000011011;
12'd950 : tab = 23'b00111101010110101010100;
12'd951 : tab = 23'b00111101010011010010000;
12'd952 : tab = 23'b00111101001111111001011;
12'd953 : tab = 23'b00111101001100100000111;
12'd954 : tab = 23'b00111101001001001000100;
12'd955 : tab = 23'b00111101000101110000001;
12'd956 : tab = 23'b00111101000010011000000;
12'd957 : tab = 23'b00111100111111000000000;
12'd958 : tab = 23'b00111100111011101000000;
12'd959 : tab = 23'b00111100111000010000010;
12'd960 : tab = 23'b00111100110100111000011;
12'd961 : tab = 23'b00111100110001100000111;
12'd962 : tab = 23'b00111100101110001001011;
12'd963 : tab = 23'b00111100101010110001111;
12'd964 : tab = 23'b00111100100111011010100;
12'd965 : tab = 23'b00111100100100000011100;
12'd966 : tab = 23'b00111100100000101100011;
12'd967 : tab = 23'b00111100011101010101011;
12'd968 : tab = 23'b00111100011001111110100;
12'd969 : tab = 23'b00111100010110100111110;
12'd970 : tab = 23'b00111100010011010001001;
12'd971 : tab = 23'b00111100001111111010101;
12'd972 : tab = 23'b00111100001100100100000;
12'd973 : tab = 23'b00111100001001001101110;
12'd974 : tab = 23'b00111100000101110111100;
12'd975 : tab = 23'b00111100000010100001011;
12'd976 : tab = 23'b00111011111111001011011;
12'd977 : tab = 23'b00111011111011110101100;
12'd978 : tab = 23'b00111011111000011111101;
12'd979 : tab = 23'b00111011110101001001111;
12'd980 : tab = 23'b00111011110001110100011;
12'd981 : tab = 23'b00111011101110011110111;
12'd982 : tab = 23'b00111011101011001001100;
12'd983 : tab = 23'b00111011100111110100001;
12'd984 : tab = 23'b00111011100100011111000;
12'd985 : tab = 23'b00111011100001001010000;
12'd986 : tab = 23'b00111011011101110101000;
12'd987 : tab = 23'b00111011011010100000001;
12'd988 : tab = 23'b00111011010111001011010;
12'd989 : tab = 23'b00111011010011110110110;
12'd990 : tab = 23'b00111011010000100010010;
12'd991 : tab = 23'b00111011001101001101110;
12'd992 : tab = 23'b00111011001001111001011;
12'd993 : tab = 23'b00111011000110100101010;
12'd994 : tab = 23'b00111011000011010001000;
12'd995 : tab = 23'b00111010111111111101000;
12'd996 : tab = 23'b00111010111100101001001;
12'd997 : tab = 23'b00111010111001010101011;
12'd998 : tab = 23'b00111010110110000001101;
12'd999 : tab = 23'b00111010110010101110000;
12'd1000 : tab = 23'b00111010101111011010100;
12'd1001 : tab = 23'b00111010101100000111001;
12'd1002 : tab = 23'b00111010101000110100000;
12'd1003 : tab = 23'b00111010100101100000101;
12'd1004 : tab = 23'b00111010100010001101101;
12'd1005 : tab = 23'b00111010011110111010100;
12'd1006 : tab = 23'b00111010011011100111101;
12'd1007 : tab = 23'b00111010011000010101000;
12'd1008 : tab = 23'b00111010010101000010010;
12'd1009 : tab = 23'b00111010010001101111110;
12'd1010 : tab = 23'b00111010001110011101010;
12'd1011 : tab = 23'b00111010001011001011000;
12'd1012 : tab = 23'b00111010000111111000101;
12'd1013 : tab = 23'b00111010000100100110100;
12'd1014 : tab = 23'b00111010000001010100100;
12'd1015 : tab = 23'b00111001111110000010100;
12'd1016 : tab = 23'b00111001111010110000110;
12'd1017 : tab = 23'b00111001110111011110111;
12'd1018 : tab = 23'b00111001110100001101010;
12'd1019 : tab = 23'b00111001110000111011110;
12'd1020 : tab = 23'b00111001101101101010010;
12'd1021 : tab = 23'b00111001101010011001000;
12'd1022 : tab = 23'b00111001100111000111110;
12'd1023 : tab = 23'b00111001100011110110101;
12'd1024 : tab = 23'b00111001100000100101101;
12'd1025 : tab = 23'b00111001011101010100101;
12'd1026 : tab = 23'b00111001011010000100000;
12'd1027 : tab = 23'b00111001010110110011001;
12'd1028 : tab = 23'b00111001010011100010100;
12'd1029 : tab = 23'b00111001010000010010000;
12'd1030 : tab = 23'b00111001001101000001100;
12'd1031 : tab = 23'b00111001001001110001010;
12'd1032 : tab = 23'b00111001000110100001001;
12'd1033 : tab = 23'b00111001000011010001000;
12'd1034 : tab = 23'b00111001000000000001000;
12'd1035 : tab = 23'b00111000111100110001001;
12'd1036 : tab = 23'b00111000111001100001010;
12'd1037 : tab = 23'b00111000110110010001101;
12'd1038 : tab = 23'b00111000110011000010000;
12'd1039 : tab = 23'b00111000101111110010100;
12'd1040 : tab = 23'b00111000101100100011001;
12'd1041 : tab = 23'b00111000101001010011110;
12'd1042 : tab = 23'b00111000100110000100100;
12'd1043 : tab = 23'b00111000100010110101100;
12'd1044 : tab = 23'b00111000011111100110100;
12'd1045 : tab = 23'b00111000011100010111100;
12'd1046 : tab = 23'b00111000011001001000110;
12'd1047 : tab = 23'b00111000010101111010001;
12'd1048 : tab = 23'b00111000010010101011100;
12'd1049 : tab = 23'b00111000001111011101000;
12'd1050 : tab = 23'b00111000001100001110101;
12'd1051 : tab = 23'b00111000001001000000011;
12'd1052 : tab = 23'b00111000000101110010000;
12'd1053 : tab = 23'b00111000000010100100000;
12'd1054 : tab = 23'b00110111111111010110000;
12'd1055 : tab = 23'b00110111111100001000001;
12'd1056 : tab = 23'b00110111111000111010010;
12'd1057 : tab = 23'b00110111110101101100100;
12'd1058 : tab = 23'b00110111110010011111000;
12'd1059 : tab = 23'b00110111101111010001100;
12'd1060 : tab = 23'b00110111101100000100000;
12'd1061 : tab = 23'b00110111101000110110110;
12'd1062 : tab = 23'b00110111100101101001101;
12'd1063 : tab = 23'b00110111100010011100100;
12'd1064 : tab = 23'b00110111011111001111011;
12'd1065 : tab = 23'b00110111011100000010100;
12'd1066 : tab = 23'b00110111011000110101110;
12'd1067 : tab = 23'b00110111010101101001000;
12'd1068 : tab = 23'b00110111010010011100100;
12'd1069 : tab = 23'b00110111001111010000000;
12'd1070 : tab = 23'b00110111001100000011100;
12'd1071 : tab = 23'b00110111001000110111010;
12'd1072 : tab = 23'b00110111000101101011000;
12'd1073 : tab = 23'b00110111000010011110111;
12'd1074 : tab = 23'b00110110111111010010111;
12'd1075 : tab = 23'b00110110111100000110111;
12'd1076 : tab = 23'b00110110111000111011000;
12'd1077 : tab = 23'b00110110110101101111100;
12'd1078 : tab = 23'b00110110110010100011110;
12'd1079 : tab = 23'b00110110101111011000010;
12'd1080 : tab = 23'b00110110101100001100110;
12'd1081 : tab = 23'b00110110101001000001100;
12'd1082 : tab = 23'b00110110100101110110001;
12'd1083 : tab = 23'b00110110100010101011001;
12'd1084 : tab = 23'b00110110011111100000000;
12'd1085 : tab = 23'b00110110011100010101000;
12'd1086 : tab = 23'b00110110011001001010010;
12'd1087 : tab = 23'b00110110010101111111100;
12'd1088 : tab = 23'b00110110010010110100110;
12'd1089 : tab = 23'b00110110001111101010001;
12'd1090 : tab = 23'b00110110001100011111110;
12'd1091 : tab = 23'b00110110001001010101011;
12'd1092 : tab = 23'b00110110000110001011001;
12'd1093 : tab = 23'b00110110000011000000111;
12'd1094 : tab = 23'b00110101111111110111000;
12'd1095 : tab = 23'b00110101111100101100110;
12'd1096 : tab = 23'b00110101111001100011000;
12'd1097 : tab = 23'b00110101110110011001010;
12'd1098 : tab = 23'b00110101110011001111100;
12'd1099 : tab = 23'b00110101110000000101111;
12'd1100 : tab = 23'b00110101101100111100100;
12'd1101 : tab = 23'b00110101101001110011000;
12'd1102 : tab = 23'b00110101100110101001110;
12'd1103 : tab = 23'b00110101100011100000100;
12'd1104 : tab = 23'b00110101100000010111010;
12'd1105 : tab = 23'b00110101011101001110011;
12'd1106 : tab = 23'b00110101011010000101011;
12'd1107 : tab = 23'b00110101010110111100110;
12'd1108 : tab = 23'b00110101010011110011111;
12'd1109 : tab = 23'b00110101010000101011010;
12'd1110 : tab = 23'b00110101001101100010101;
12'd1111 : tab = 23'b00110101001010011010010;
12'd1112 : tab = 23'b00110101000111010010000;
12'd1113 : tab = 23'b00110101000100001001110;
12'd1114 : tab = 23'b00110101000001000001100;
12'd1115 : tab = 23'b00110100111101111001011;
12'd1116 : tab = 23'b00110100111010110001011;
12'd1117 : tab = 23'b00110100110111101001101;
12'd1118 : tab = 23'b00110100110100100001110;
12'd1119 : tab = 23'b00110100110001011010000;
12'd1120 : tab = 23'b00110100101110010010100;
12'd1121 : tab = 23'b00110100101011001011000;
12'd1122 : tab = 23'b00110100101000000011100;
12'd1123 : tab = 23'b00110100100100111100010;
12'd1124 : tab = 23'b00110100100001110101000;
12'd1125 : tab = 23'b00110100011110101110000;
12'd1126 : tab = 23'b00110100011011100110111;
12'd1127 : tab = 23'b00110100011000100000000;
12'd1128 : tab = 23'b00110100010101011001010;
12'd1129 : tab = 23'b00110100010010010010011;
12'd1130 : tab = 23'b00110100001111001011110;
12'd1131 : tab = 23'b00110100001100000101001;
12'd1132 : tab = 23'b00110100001000111110101;
12'd1133 : tab = 23'b00110100000101111000011;
12'd1134 : tab = 23'b00110100000010110010000;
12'd1135 : tab = 23'b00110011111111101011111;
12'd1136 : tab = 23'b00110011111100100101110;
12'd1137 : tab = 23'b00110011111001011111110;
12'd1138 : tab = 23'b00110011110110011001110;
12'd1139 : tab = 23'b00110011110011010100001;
12'd1140 : tab = 23'b00110011110000001110010;
12'd1141 : tab = 23'b00110011101101001000110;
12'd1142 : tab = 23'b00110011101010000011001;
12'd1143 : tab = 23'b00110011100110111101110;
12'd1144 : tab = 23'b00110011100011111000011;
12'd1145 : tab = 23'b00110011100000110011001;
12'd1146 : tab = 23'b00110011011101101110000;
12'd1147 : tab = 23'b00110011011010101000111;
12'd1148 : tab = 23'b00110011010111100100000;
12'd1149 : tab = 23'b00110011010100011111000;
12'd1150 : tab = 23'b00110011010001011010010;
12'd1151 : tab = 23'b00110011001110010101100;
12'd1152 : tab = 23'b00110011001011010000111;
12'd1153 : tab = 23'b00110011001000001100011;
12'd1154 : tab = 23'b00110011000101001000000;
12'd1155 : tab = 23'b00110011000010000011110;
12'd1156 : tab = 23'b00110010111110111111100;
12'd1157 : tab = 23'b00110010111011111011010;
12'd1158 : tab = 23'b00110010111000110111010;
12'd1159 : tab = 23'b00110010110101110011010;
12'd1160 : tab = 23'b00110010110010101111010;
12'd1161 : tab = 23'b00110010101111101011100;
12'd1162 : tab = 23'b00110010101100100111111;
12'd1163 : tab = 23'b00110010101001100100010;
12'd1164 : tab = 23'b00110010100110100000111;
12'd1165 : tab = 23'b00110010100011011101010;
12'd1166 : tab = 23'b00110010100000011010000;
12'd1167 : tab = 23'b00110010011101010111000;
12'd1168 : tab = 23'b00110010011010010011101;
12'd1169 : tab = 23'b00110010010111010000110;
12'd1170 : tab = 23'b00110010010100001101101;
12'd1171 : tab = 23'b00110010010001001010110;
12'd1172 : tab = 23'b00110010001110001000000;
12'd1173 : tab = 23'b00110010001011000101010;
12'd1174 : tab = 23'b00110010001000000010110;
12'd1175 : tab = 23'b00110010000101000000010;
12'd1176 : tab = 23'b00110010000001111101110;
12'd1177 : tab = 23'b00110001111110111011100;
12'd1178 : tab = 23'b00110001111011111001010;
12'd1179 : tab = 23'b00110001111000110111000;
12'd1180 : tab = 23'b00110001110101110101000;
12'd1181 : tab = 23'b00110001110010110011001;
12'd1182 : tab = 23'b00110001101111110001010;
12'd1183 : tab = 23'b00110001101100101111100;
12'd1184 : tab = 23'b00110001101001101101110;
12'd1185 : tab = 23'b00110001100110101100001;
12'd1186 : tab = 23'b00110001100011101010101;
12'd1187 : tab = 23'b00110001100000101001010;
12'd1188 : tab = 23'b00110001011101100111111;
12'd1189 : tab = 23'b00110001011010100110100;
12'd1190 : tab = 23'b00110001010111100101100;
12'd1191 : tab = 23'b00110001010100100100011;
12'd1192 : tab = 23'b00110001010001100011100;
12'd1193 : tab = 23'b00110001001110100010100;
12'd1194 : tab = 23'b00110001001011100001110;
12'd1195 : tab = 23'b00110001001000100001000;
12'd1196 : tab = 23'b00110001000101100000100;
12'd1197 : tab = 23'b00110001000010011111110;
12'd1198 : tab = 23'b00110000111111011111100;
12'd1199 : tab = 23'b00110000111100011111000;
12'd1200 : tab = 23'b00110000111001011110111;
12'd1201 : tab = 23'b00110000110110011110101;
12'd1202 : tab = 23'b00110000110011011110100;
12'd1203 : tab = 23'b00110000110000011110100;
12'd1204 : tab = 23'b00110000101101011110110;
12'd1205 : tab = 23'b00110000101010011110110;
12'd1206 : tab = 23'b00110000100111011111000;
12'd1207 : tab = 23'b00110000100100011111100;
12'd1208 : tab = 23'b00110000100001011111110;
12'd1209 : tab = 23'b00110000011110100000011;
12'd1210 : tab = 23'b00110000011011100001000;
12'd1211 : tab = 23'b00110000011000100001110;
12'd1212 : tab = 23'b00110000010101100010101;
12'd1213 : tab = 23'b00110000010010100011011;
12'd1214 : tab = 23'b00110000001111100100010;
12'd1215 : tab = 23'b00110000001100100101100;
12'd1216 : tab = 23'b00110000001001100110100;
12'd1217 : tab = 23'b00110000000110100111110;
12'd1218 : tab = 23'b00110000000011101001000;
12'd1219 : tab = 23'b00110000000000101010100;
12'd1220 : tab = 23'b00101111111101101100000;
12'd1221 : tab = 23'b00101111111010101101101;
12'd1222 : tab = 23'b00101111110111101111010;
12'd1223 : tab = 23'b00101111110100110001000;
12'd1224 : tab = 23'b00101111110001110011000;
12'd1225 : tab = 23'b00101111101110110100110;
12'd1226 : tab = 23'b00101111101011110110111;
12'd1227 : tab = 23'b00101111101000111001000;
12'd1228 : tab = 23'b00101111100101111011010;
12'd1229 : tab = 23'b00101111100010111101100;
12'd1230 : tab = 23'b00101111011111111111110;
12'd1231 : tab = 23'b00101111011101000010010;
12'd1232 : tab = 23'b00101111011010000100110;
12'd1233 : tab = 23'b00101111010111000111011;
12'd1234 : tab = 23'b00101111010100001010010;
12'd1235 : tab = 23'b00101111010001001100110;
12'd1236 : tab = 23'b00101111001110001111110;
12'd1237 : tab = 23'b00101111001011010010110;
12'd1238 : tab = 23'b00101111001000010101110;
12'd1239 : tab = 23'b00101111000101011001000;
12'd1240 : tab = 23'b00101111000010011100010;
12'd1241 : tab = 23'b00101110111111011111100;
12'd1242 : tab = 23'b00101110111100100011000;
12'd1243 : tab = 23'b00101110111001100110100;
12'd1244 : tab = 23'b00101110110110101001111;
12'd1245 : tab = 23'b00101110110011101101101;
12'd1246 : tab = 23'b00101110110000110001011;
12'd1247 : tab = 23'b00101110101101110101010;
12'd1248 : tab = 23'b00101110101010111001001;
12'd1249 : tab = 23'b00101110100111111101010;
12'd1250 : tab = 23'b00101110100101000001010;
12'd1251 : tab = 23'b00101110100010000101100;
12'd1252 : tab = 23'b00101110011111001001110;
12'd1253 : tab = 23'b00101110011100001110000;
12'd1254 : tab = 23'b00101110011001010010100;
12'd1255 : tab = 23'b00101110010110010111000;
12'd1256 : tab = 23'b00101110010011011011100;
12'd1257 : tab = 23'b00101110010000100000010;
12'd1258 : tab = 23'b00101110001101100101000;
12'd1259 : tab = 23'b00101110001010101010000;
12'd1260 : tab = 23'b00101110000111101110111;
12'd1261 : tab = 23'b00101110000100110011111;
12'd1262 : tab = 23'b00101110000001111001000;
12'd1263 : tab = 23'b00101101111110111110010;
12'd1264 : tab = 23'b00101101111100000011011;
12'd1265 : tab = 23'b00101101111001001000110;
12'd1266 : tab = 23'b00101101110110001110010;
12'd1267 : tab = 23'b00101101110011010011110;
12'd1268 : tab = 23'b00101101110000011001100;
12'd1269 : tab = 23'b00101101101101011111000;
12'd1270 : tab = 23'b00101101101010100100111;
12'd1271 : tab = 23'b00101101100111101010110;
12'd1272 : tab = 23'b00101101100100110000110;
12'd1273 : tab = 23'b00101101100001110110110;
12'd1274 : tab = 23'b00101101011110111100111;
12'd1275 : tab = 23'b00101101011100000011000;
12'd1276 : tab = 23'b00101101011001001001011;
12'd1277 : tab = 23'b00101101010110001111110;
12'd1278 : tab = 23'b00101101010011010110010;
12'd1279 : tab = 23'b00101101010000011100110;
12'd1280 : tab = 23'b00101101001101100011011;
12'd1281 : tab = 23'b00101101001010101010001;
12'd1282 : tab = 23'b00101101000111110000111;
12'd1283 : tab = 23'b00101101000100110111110;
12'd1284 : tab = 23'b00101101000001111110110;
12'd1285 : tab = 23'b00101100111111000101110;
12'd1286 : tab = 23'b00101100111100001101000;
12'd1287 : tab = 23'b00101100111001010100000;
12'd1288 : tab = 23'b00101100110110011011011;
12'd1289 : tab = 23'b00101100110011100010111;
12'd1290 : tab = 23'b00101100110000101010010;
12'd1291 : tab = 23'b00101100101101110001110;
12'd1292 : tab = 23'b00101100101010111001011;
12'd1293 : tab = 23'b00101100101000000001000;
12'd1294 : tab = 23'b00101100100101001001000;
12'd1295 : tab = 23'b00101100100010010000110;
12'd1296 : tab = 23'b00101100011111011000110;
12'd1297 : tab = 23'b00101100011100100000110;
12'd1298 : tab = 23'b00101100011001101000111;
12'd1299 : tab = 23'b00101100010110110001000;
12'd1300 : tab = 23'b00101100010011111001010;
12'd1301 : tab = 23'b00101100010001000001110;
12'd1302 : tab = 23'b00101100001110001010010;
12'd1303 : tab = 23'b00101100001011010010101;
12'd1304 : tab = 23'b00101100001000011011010;
12'd1305 : tab = 23'b00101100000101100100000;
12'd1306 : tab = 23'b00101100000010101100110;
12'd1307 : tab = 23'b00101011111111110101110;
12'd1308 : tab = 23'b00101011111100111110101;
12'd1309 : tab = 23'b00101011111010000111101;
12'd1310 : tab = 23'b00101011110111010000110;
12'd1311 : tab = 23'b00101011110100011001111;
12'd1312 : tab = 23'b00101011110001100011001;
12'd1313 : tab = 23'b00101011101110101100100;
12'd1314 : tab = 23'b00101011101011110101111;
12'd1315 : tab = 23'b00101011101000111111100;
12'd1316 : tab = 23'b00101011100110001001000;
12'd1317 : tab = 23'b00101011100011010010110;
12'd1318 : tab = 23'b00101011100000011100100;
12'd1319 : tab = 23'b00101011011101100110011;
12'd1320 : tab = 23'b00101011011010110000010;
12'd1321 : tab = 23'b00101011010111111010010;
12'd1322 : tab = 23'b00101011010101000100010;
12'd1323 : tab = 23'b00101011010010001110100;
12'd1324 : tab = 23'b00101011001111011000101;
12'd1325 : tab = 23'b00101011001100100011000;
12'd1326 : tab = 23'b00101011001001101101100;
12'd1327 : tab = 23'b00101011000110110111111;
12'd1328 : tab = 23'b00101011000100000010100;
12'd1329 : tab = 23'b00101011000001001101001;
12'd1330 : tab = 23'b00101010111110010111110;
12'd1331 : tab = 23'b00101010111011100010110;
12'd1332 : tab = 23'b00101010111000101101100;
12'd1333 : tab = 23'b00101010110101111000100;
12'd1334 : tab = 23'b00101010110011000011100;
12'd1335 : tab = 23'b00101010110000001110101;
12'd1336 : tab = 23'b00101010101101011001111;
12'd1337 : tab = 23'b00101010101010100101010;
12'd1338 : tab = 23'b00101010100111110000100;
12'd1339 : tab = 23'b00101010100100111100000;
12'd1340 : tab = 23'b00101010100010000111100;
12'd1341 : tab = 23'b00101010011111010011001;
12'd1342 : tab = 23'b00101010011100011110110;
12'd1343 : tab = 23'b00101010011001101010101;
12'd1344 : tab = 23'b00101010010110110110100;
12'd1345 : tab = 23'b00101010010100000010010;
12'd1346 : tab = 23'b00101010010001001110011;
12'd1347 : tab = 23'b00101010001110011010100;
12'd1348 : tab = 23'b00101010001011100110101;
12'd1349 : tab = 23'b00101010001000110010110;
12'd1350 : tab = 23'b00101010000101111111010;
12'd1351 : tab = 23'b00101010000011001011100;
12'd1352 : tab = 23'b00101010000000011000000;
12'd1353 : tab = 23'b00101001111101100100110;
12'd1354 : tab = 23'b00101001111010110001010;
12'd1355 : tab = 23'b00101001110111111110000;
12'd1356 : tab = 23'b00101001110101001010110;
12'd1357 : tab = 23'b00101001110010010111110;
12'd1358 : tab = 23'b00101001101111100100101;
12'd1359 : tab = 23'b00101001101100110001100;
12'd1360 : tab = 23'b00101001101001111110110;
12'd1361 : tab = 23'b00101001100111001100000;
12'd1362 : tab = 23'b00101001100100011001010;
12'd1363 : tab = 23'b00101001100001100110101;
12'd1364 : tab = 23'b00101001011110110100000;
12'd1365 : tab = 23'b00101001011100000001100;
12'd1366 : tab = 23'b00101001011001001111001;
12'd1367 : tab = 23'b00101001010110011100110;
12'd1368 : tab = 23'b00101001010011101010100;
12'd1369 : tab = 23'b00101001010000111000010;
12'd1370 : tab = 23'b00101001001110000110010;
12'd1371 : tab = 23'b00101001001011010100001;
12'd1372 : tab = 23'b00101001001000100010010;
12'd1373 : tab = 23'b00101001000101110000011;
12'd1374 : tab = 23'b00101001000010111110101;
12'd1375 : tab = 23'b00101001000000001101000;
12'd1376 : tab = 23'b00101000111101011011010;
12'd1377 : tab = 23'b00101000111010101001110;
12'd1378 : tab = 23'b00101000110111111000001;
12'd1379 : tab = 23'b00101000110101000110110;
12'd1380 : tab = 23'b00101000110010010101100;
12'd1381 : tab = 23'b00101000101111100100010;
12'd1382 : tab = 23'b00101000101100110011001;
12'd1383 : tab = 23'b00101000101010000010000;
12'd1384 : tab = 23'b00101000100111010001000;
12'd1385 : tab = 23'b00101000100100100000000;
12'd1386 : tab = 23'b00101000100001101111001;
12'd1387 : tab = 23'b00101000011110111110100;
12'd1388 : tab = 23'b00101000011100001101110;
12'd1389 : tab = 23'b00101000011001011101000;
12'd1390 : tab = 23'b00101000010110101100100;
12'd1391 : tab = 23'b00101000010011111100000;
12'd1392 : tab = 23'b00101000010001001011110;
12'd1393 : tab = 23'b00101000001110011011010;
12'd1394 : tab = 23'b00101000001011101011000;
12'd1395 : tab = 23'b00101000001000111010111;
12'd1396 : tab = 23'b00101000000110001010111;
12'd1397 : tab = 23'b00101000000011011010110;
12'd1398 : tab = 23'b00101000000000101010110;
12'd1399 : tab = 23'b00100111111101111011001;
12'd1400 : tab = 23'b00100111111011001011010;
12'd1401 : tab = 23'b00100111111000011011100;
12'd1402 : tab = 23'b00100111110101101100000;
12'd1403 : tab = 23'b00100111110010111100011;
12'd1404 : tab = 23'b00100111110000001100111;
12'd1405 : tab = 23'b00100111101101011101011;
12'd1406 : tab = 23'b00100111101010101110001;
12'd1407 : tab = 23'b00100111100111111111000;
12'd1408 : tab = 23'b00100111100101001111110;
12'd1409 : tab = 23'b00100111100010100000110;
12'd1410 : tab = 23'b00100111011111110001100;
12'd1411 : tab = 23'b00100111011101000010101;
12'd1412 : tab = 23'b00100111011010010011110;
12'd1413 : tab = 23'b00100111010111100101000;
12'd1414 : tab = 23'b00100111010100110110010;
12'd1415 : tab = 23'b00100111010010000111101;
12'd1416 : tab = 23'b00100111001111011001000;
12'd1417 : tab = 23'b00100111001100101010101;
12'd1418 : tab = 23'b00100111001001111100001;
12'd1419 : tab = 23'b00100111000111001101111;
12'd1420 : tab = 23'b00100111000100011111100;
12'd1421 : tab = 23'b00100111000001110001011;
12'd1422 : tab = 23'b00100110111111000011010;
12'd1423 : tab = 23'b00100110111100010101010;
12'd1424 : tab = 23'b00100110111001100111010;
12'd1425 : tab = 23'b00100110110110111001011;
12'd1426 : tab = 23'b00100110110100001011100;
12'd1427 : tab = 23'b00100110110001011101110;
12'd1428 : tab = 23'b00100110101110110000001;
12'd1429 : tab = 23'b00100110101100000010101;
12'd1430 : tab = 23'b00100110101001010101000;
12'd1431 : tab = 23'b00100110100110100111101;
12'd1432 : tab = 23'b00100110100011111010010;
12'd1433 : tab = 23'b00100110100001001101000;
12'd1434 : tab = 23'b00100110011110011111110;
12'd1435 : tab = 23'b00100110011011110010101;
12'd1436 : tab = 23'b00100110011001000101100;
12'd1437 : tab = 23'b00100110010110011000101;
12'd1438 : tab = 23'b00100110010011101011101;
12'd1439 : tab = 23'b00100110010000111111000;
12'd1440 : tab = 23'b00100110001110010010000;
12'd1441 : tab = 23'b00100110001011100101011;
12'd1442 : tab = 23'b00100110001000111000110;
12'd1443 : tab = 23'b00100110000110001100010;
12'd1444 : tab = 23'b00100110000011011111110;
12'd1445 : tab = 23'b00100110000000110011011;
12'd1446 : tab = 23'b00100101111110000111000;
12'd1447 : tab = 23'b00100101111011011010110;
12'd1448 : tab = 23'b00100101111000101110101;
12'd1449 : tab = 23'b00100101110110000010100;
12'd1450 : tab = 23'b00100101110011010110011;
12'd1451 : tab = 23'b00100101110000101010100;
12'd1452 : tab = 23'b00100101101101111110110;
12'd1453 : tab = 23'b00100101101011010010110;
12'd1454 : tab = 23'b00100101101000100111000;
12'd1455 : tab = 23'b00100101100101111011100;
12'd1456 : tab = 23'b00100101100011001111111;
12'd1457 : tab = 23'b00100101100000100100010;
12'd1458 : tab = 23'b00100101011101111000111;
12'd1459 : tab = 23'b00100101011011001101100;
12'd1460 : tab = 23'b00100101011000100010010;
12'd1461 : tab = 23'b00100101010101110111000;
12'd1462 : tab = 23'b00100101010011001011110;
12'd1463 : tab = 23'b00100101010000100000110;
12'd1464 : tab = 23'b00100101001101110101110;
12'd1465 : tab = 23'b00100101001011001010110;
12'd1466 : tab = 23'b00100101001000100000000;
12'd1467 : tab = 23'b00100101000101110101010;
12'd1468 : tab = 23'b00100101000011001010100;
12'd1469 : tab = 23'b00100101000000100000000;
12'd1470 : tab = 23'b00100100111101110101010;
12'd1471 : tab = 23'b00100100111011001010111;
12'd1472 : tab = 23'b00100100111000100000100;
12'd1473 : tab = 23'b00100100110101110110001;
12'd1474 : tab = 23'b00100100110011001011110;
12'd1475 : tab = 23'b00100100110000100001110;
12'd1476 : tab = 23'b00100100101101110111100;
12'd1477 : tab = 23'b00100100101011001101011;
12'd1478 : tab = 23'b00100100101000100011011;
12'd1479 : tab = 23'b00100100100101111001100;
12'd1480 : tab = 23'b00100100100011001111110;
12'd1481 : tab = 23'b00100100100000100101111;
12'd1482 : tab = 23'b00100100011101111100010;
12'd1483 : tab = 23'b00100100011011010010110;
12'd1484 : tab = 23'b00100100011000101001000;
12'd1485 : tab = 23'b00100100010101111111101;
12'd1486 : tab = 23'b00100100010011010110010;
12'd1487 : tab = 23'b00100100010000101100111;
12'd1488 : tab = 23'b00100100001110000011100;
12'd1489 : tab = 23'b00100100001011011010100;
12'd1490 : tab = 23'b00100100001000110001010;
12'd1491 : tab = 23'b00100100000110001000010;
12'd1492 : tab = 23'b00100100000011011111010;
12'd1493 : tab = 23'b00100100000000110110010;
12'd1494 : tab = 23'b00100011111110001101100;
12'd1495 : tab = 23'b00100011111011100100110;
12'd1496 : tab = 23'b00100011111000111100000;
12'd1497 : tab = 23'b00100011110110010011011;
12'd1498 : tab = 23'b00100011110011101011000;
12'd1499 : tab = 23'b00100011110001000010100;
12'd1500 : tab = 23'b00100011101110011010000;
12'd1501 : tab = 23'b00100011101011110001110;
12'd1502 : tab = 23'b00100011101001001001100;
12'd1503 : tab = 23'b00100011100110100001010;
12'd1504 : tab = 23'b00100011100011111001001;
12'd1505 : tab = 23'b00100011100001010001000;
12'd1506 : tab = 23'b00100011011110101001000;
12'd1507 : tab = 23'b00100011011100000001010;
12'd1508 : tab = 23'b00100011011001011001100;
12'd1509 : tab = 23'b00100011010110110001101;
12'd1510 : tab = 23'b00100011010100001001111;
12'd1511 : tab = 23'b00100011010001100010011;
12'd1512 : tab = 23'b00100011001110111010110;
12'd1513 : tab = 23'b00100011001100010011010;
12'd1514 : tab = 23'b00100011001001101011111;
12'd1515 : tab = 23'b00100011000111000100100;
12'd1516 : tab = 23'b00100011000100011101010;
12'd1517 : tab = 23'b00100011000001110110000;
12'd1518 : tab = 23'b00100010111111001110111;
12'd1519 : tab = 23'b00100010111100100111110;
12'd1520 : tab = 23'b00100010111010000001000;
12'd1521 : tab = 23'b00100010110111011001111;
12'd1522 : tab = 23'b00100010110100110011000;
12'd1523 : tab = 23'b00100010110010001100010;
12'd1524 : tab = 23'b00100010101111100101101;
12'd1525 : tab = 23'b00100010101100111111000;
12'd1526 : tab = 23'b00100010101010011000011;
12'd1527 : tab = 23'b00100010100111110010000;
12'd1528 : tab = 23'b00100010100101001011100;
12'd1529 : tab = 23'b00100010100010100101001;
12'd1530 : tab = 23'b00100010011111111110110;
12'd1531 : tab = 23'b00100010011101011000100;
12'd1532 : tab = 23'b00100010011010110010011;
12'd1533 : tab = 23'b00100010011000001100011;
12'd1534 : tab = 23'b00100010010101100110010;
12'd1535 : tab = 23'b00100010010011000000011;
12'd1536 : tab = 23'b00100010010000011010101;
12'd1537 : tab = 23'b00100010001101110100110;
12'd1538 : tab = 23'b00100010001011001111000;
12'd1539 : tab = 23'b00100010001000101001010;
12'd1540 : tab = 23'b00100010000110000011110;
12'd1541 : tab = 23'b00100010000011011110010;
12'd1542 : tab = 23'b00100010000000111000110;
12'd1543 : tab = 23'b00100001111110010011010;
12'd1544 : tab = 23'b00100001111011101110000;
12'd1545 : tab = 23'b00100001111001001000110;
12'd1546 : tab = 23'b00100001110110100011100;
12'd1547 : tab = 23'b00100001110011111110100;
12'd1548 : tab = 23'b00100001110001011001100;
12'd1549 : tab = 23'b00100001101110110100100;
12'd1550 : tab = 23'b00100001101100001111100;
12'd1551 : tab = 23'b00100001101001101010110;
12'd1552 : tab = 23'b00100001100111000110000;
12'd1553 : tab = 23'b00100001100100100001010;
12'd1554 : tab = 23'b00100001100001111100110;
12'd1555 : tab = 23'b00100001011111011000000;
12'd1556 : tab = 23'b00100001011100110011101;
12'd1557 : tab = 23'b00100001011010001111010;
12'd1558 : tab = 23'b00100001010111101010111;
12'd1559 : tab = 23'b00100001010101000110100;
12'd1560 : tab = 23'b00100001010010100010010;
12'd1561 : tab = 23'b00100001001111111110001;
12'd1562 : tab = 23'b00100001001101011010001;
12'd1563 : tab = 23'b00100001001010110110000;
12'd1564 : tab = 23'b00100001001000010010001;
12'd1565 : tab = 23'b00100001000101101110010;
12'd1566 : tab = 23'b00100001000011001010100;
12'd1567 : tab = 23'b00100001000000100110110;
12'd1568 : tab = 23'b00100000111110000011000;
12'd1569 : tab = 23'b00100000111011011111011;
12'd1570 : tab = 23'b00100000111000111011111;
12'd1571 : tab = 23'b00100000110110011000011;
12'd1572 : tab = 23'b00100000110011110101000;
12'd1573 : tab = 23'b00100000110001010001101;
12'd1574 : tab = 23'b00100000101110101110011;
12'd1575 : tab = 23'b00100000101100001011001;
12'd1576 : tab = 23'b00100000101001101000000;
12'd1577 : tab = 23'b00100000100111000100111;
12'd1578 : tab = 23'b00100000100100100010000;
12'd1579 : tab = 23'b00100000100001111111000;
12'd1580 : tab = 23'b00100000011111011100001;
12'd1581 : tab = 23'b00100000011100111001011;
12'd1582 : tab = 23'b00100000011010010110100;
12'd1583 : tab = 23'b00100000010111110100000;
12'd1584 : tab = 23'b00100000010101010001100;
12'd1585 : tab = 23'b00100000010010101110111;
12'd1586 : tab = 23'b00100000010000001100011;
12'd1587 : tab = 23'b00100000001101101010000;
12'd1588 : tab = 23'b00100000001011000111101;
12'd1589 : tab = 23'b00100000001000100101011;
12'd1590 : tab = 23'b00100000000110000011010;
12'd1591 : tab = 23'b00100000000011100001001;
12'd1592 : tab = 23'b00100000000000111111000;
12'd1593 : tab = 23'b00011111111110011101000;
12'd1594 : tab = 23'b00011111111011111011010;
12'd1595 : tab = 23'b00011111111001011001010;
12'd1596 : tab = 23'b00011111110110110111100;
12'd1597 : tab = 23'b00011111110100010101110;
12'd1598 : tab = 23'b00011111110001110100001;
12'd1599 : tab = 23'b00011111101111010010100;
12'd1600 : tab = 23'b00011111101100110001000;
12'd1601 : tab = 23'b00011111101010001111100;
12'd1602 : tab = 23'b00011111100111101110001;
12'd1603 : tab = 23'b00011111100101001100110;
12'd1604 : tab = 23'b00011111100010101011100;
12'd1605 : tab = 23'b00011111100000001010010;
12'd1606 : tab = 23'b00011111011101101001010;
12'd1607 : tab = 23'b00011111011011001000001;
12'd1608 : tab = 23'b00011111011000100111000;
12'd1609 : tab = 23'b00011111010110000110010;
12'd1610 : tab = 23'b00011111010011100101010;
12'd1611 : tab = 23'b00011111010001000100100;
12'd1612 : tab = 23'b00011111001110100011110;
12'd1613 : tab = 23'b00011111001100000011000;
12'd1614 : tab = 23'b00011111001001100010100;
12'd1615 : tab = 23'b00011111000111000010000;
12'd1616 : tab = 23'b00011111000100100001100;
12'd1617 : tab = 23'b00011111000010000001000;
12'd1618 : tab = 23'b00011110111111100000110;
12'd1619 : tab = 23'b00011110111101000000100;
12'd1620 : tab = 23'b00011110111010100000010;
12'd1621 : tab = 23'b00011110111000000000010;
12'd1622 : tab = 23'b00011110110101100000000;
12'd1623 : tab = 23'b00011110110011000000001;
12'd1624 : tab = 23'b00011110110000100000001;
12'd1625 : tab = 23'b00011110101110000000010;
12'd1626 : tab = 23'b00011110101011100000100;
12'd1627 : tab = 23'b00011110101001000000101;
12'd1628 : tab = 23'b00011110100110100001000;
12'd1629 : tab = 23'b00011110100100000001100;
12'd1630 : tab = 23'b00011110100001100001110;
12'd1631 : tab = 23'b00011110011111000010010;
12'd1632 : tab = 23'b00011110011100100011000;
12'd1633 : tab = 23'b00011110011010000011100;
12'd1634 : tab = 23'b00011110010111100100010;
12'd1635 : tab = 23'b00011110010101000101001;
12'd1636 : tab = 23'b00011110010010100101111;
12'd1637 : tab = 23'b00011110010000000110110;
12'd1638 : tab = 23'b00011110001101100111110;
12'd1639 : tab = 23'b00011110001011001000110;
12'd1640 : tab = 23'b00011110001000101001110;
12'd1641 : tab = 23'b00011110000110001011000;
12'd1642 : tab = 23'b00011110000011101100010;
12'd1643 : tab = 23'b00011110000001001101100;
12'd1644 : tab = 23'b00011101111110101110111;
12'd1645 : tab = 23'b00011101111100010000010;
12'd1646 : tab = 23'b00011101111001110001110;
12'd1647 : tab = 23'b00011101110111010011010;
12'd1648 : tab = 23'b00011101110100110101000;
12'd1649 : tab = 23'b00011101110010010110100;
12'd1650 : tab = 23'b00011101101111111000010;
12'd1651 : tab = 23'b00011101101101011010001;
12'd1652 : tab = 23'b00011101101010111100000;
12'd1653 : tab = 23'b00011101101000011110000;
12'd1654 : tab = 23'b00011101100101111111111;
12'd1655 : tab = 23'b00011101100011100010000;
12'd1656 : tab = 23'b00011101100001000100001;
12'd1657 : tab = 23'b00011101011110100110010;
12'd1658 : tab = 23'b00011101011100001000100;
12'd1659 : tab = 23'b00011101011001101010111;
12'd1660 : tab = 23'b00011101010111001101010;
12'd1661 : tab = 23'b00011101010100101111110;
12'd1662 : tab = 23'b00011101010010010010010;
12'd1663 : tab = 23'b00011101001111110100110;
12'd1664 : tab = 23'b00011101001101010111011;
12'd1665 : tab = 23'b00011101001010111010000;
12'd1666 : tab = 23'b00011101001000011100111;
12'd1667 : tab = 23'b00011101000101111111101;
12'd1668 : tab = 23'b00011101000011100010101;
12'd1669 : tab = 23'b00011101000001000101100;
12'd1670 : tab = 23'b00011100111110101000100;
12'd1671 : tab = 23'b00011100111100001011101;
12'd1672 : tab = 23'b00011100111001101110110;
12'd1673 : tab = 23'b00011100110111010001111;
12'd1674 : tab = 23'b00011100110100110101010;
12'd1675 : tab = 23'b00011100110010011000100;
12'd1676 : tab = 23'b00011100101111111100000;
12'd1677 : tab = 23'b00011100101101011111011;
12'd1678 : tab = 23'b00011100101011000010111;
12'd1679 : tab = 23'b00011100101000100110100;
12'd1680 : tab = 23'b00011100100110001010001;
12'd1681 : tab = 23'b00011100100011101101111;
12'd1682 : tab = 23'b00011100100001010001101;
12'd1683 : tab = 23'b00011100011110110101100;
12'd1684 : tab = 23'b00011100011100011001010;
12'd1685 : tab = 23'b00011100011001111101010;
12'd1686 : tab = 23'b00011100010111100001010;
12'd1687 : tab = 23'b00011100010101000101011;
12'd1688 : tab = 23'b00011100010010101001100;
12'd1689 : tab = 23'b00011100010000001101110;
12'd1690 : tab = 23'b00011100001101110010000;
12'd1691 : tab = 23'b00011100001011010110011;
12'd1692 : tab = 23'b00011100001000111010110;
12'd1693 : tab = 23'b00011100000110011111010;
12'd1694 : tab = 23'b00011100000100000011110;
12'd1695 : tab = 23'b00011100000001101000010;
12'd1696 : tab = 23'b00011011111111001101000;
12'd1697 : tab = 23'b00011011111100110001110;
12'd1698 : tab = 23'b00011011111010010110100;
12'd1699 : tab = 23'b00011011110111111011010;
12'd1700 : tab = 23'b00011011110101100000010;
12'd1701 : tab = 23'b00011011110011000101010;
12'd1702 : tab = 23'b00011011110000101010001;
12'd1703 : tab = 23'b00011011101110001111010;
12'd1704 : tab = 23'b00011011101011110100011;
12'd1705 : tab = 23'b00011011101001011001101;
12'd1706 : tab = 23'b00011011100110111110110;
12'd1707 : tab = 23'b00011011100100100100001;
12'd1708 : tab = 23'b00011011100010001001101;
12'd1709 : tab = 23'b00011011011111101111000;
12'd1710 : tab = 23'b00011011011101010100100;
12'd1711 : tab = 23'b00011011011010111010001;
12'd1712 : tab = 23'b00011011011000011111110;
12'd1713 : tab = 23'b00011011010110000101100;
12'd1714 : tab = 23'b00011011010011101011010;
12'd1715 : tab = 23'b00011011010001010001000;
12'd1716 : tab = 23'b00011011001110110111000;
12'd1717 : tab = 23'b00011011001100011100110;
12'd1718 : tab = 23'b00011011001010000010111;
12'd1719 : tab = 23'b00011011000111101001000;
12'd1720 : tab = 23'b00011011000101001111000;
12'd1721 : tab = 23'b00011011000010110101010;
12'd1722 : tab = 23'b00011011000000011011100;
12'd1723 : tab = 23'b00011010111110000001110;
12'd1724 : tab = 23'b00011010111011101000010;
12'd1725 : tab = 23'b00011010111001001110101;
12'd1726 : tab = 23'b00011010110110110101000;
12'd1727 : tab = 23'b00011010110100011011101;
12'd1728 : tab = 23'b00011010110010000010010;
12'd1729 : tab = 23'b00011010101111101001000;
12'd1730 : tab = 23'b00011010101101001111110;
12'd1731 : tab = 23'b00011010101010110110100;
12'd1732 : tab = 23'b00011010101000011101011;
12'd1733 : tab = 23'b00011010100110000100010;
12'd1734 : tab = 23'b00011010100011101011010;
12'd1735 : tab = 23'b00011010100001010010011;
12'd1736 : tab = 23'b00011010011110111001011;
12'd1737 : tab = 23'b00011010011100100000100;
12'd1738 : tab = 23'b00011010011010000111110;
12'd1739 : tab = 23'b00011010010111101111001;
12'd1740 : tab = 23'b00011010010101010110100;
12'd1741 : tab = 23'b00011010010010111101111;
12'd1742 : tab = 23'b00011010010000100101010;
12'd1743 : tab = 23'b00011010001110001100110;
12'd1744 : tab = 23'b00011010001011110100011;
12'd1745 : tab = 23'b00011010001001011100000;
12'd1746 : tab = 23'b00011010000111000011110;
12'd1747 : tab = 23'b00011010000100101011101;
12'd1748 : tab = 23'b00011010000010010011011;
12'd1749 : tab = 23'b00011001111111111011010;
12'd1750 : tab = 23'b00011001111101100011010;
12'd1751 : tab = 23'b00011001111011001011010;
12'd1752 : tab = 23'b00011001111000110011010;
12'd1753 : tab = 23'b00011001110110011011100;
12'd1754 : tab = 23'b00011001110100000011100;
12'd1755 : tab = 23'b00011001110001101011111;
12'd1756 : tab = 23'b00011001101111010100010;
12'd1757 : tab = 23'b00011001101100111100100;
12'd1758 : tab = 23'b00011001101010100101000;
12'd1759 : tab = 23'b00011001101000001101011;
12'd1760 : tab = 23'b00011001100101110110000;
12'd1761 : tab = 23'b00011001100011011110100;
12'd1762 : tab = 23'b00011001100001000111010;
12'd1763 : tab = 23'b00011001011110110000000;
12'd1764 : tab = 23'b00011001011100011000110;
12'd1765 : tab = 23'b00011001011010000001101;
12'd1766 : tab = 23'b00011001010111101010100;
12'd1767 : tab = 23'b00011001010101010011100;
12'd1768 : tab = 23'b00011001010010111100100;
12'd1769 : tab = 23'b00011001010000100101100;
12'd1770 : tab = 23'b00011001001110001110110;
12'd1771 : tab = 23'b00011001001011110111111;
12'd1772 : tab = 23'b00011001001001100001000;
12'd1773 : tab = 23'b00011001000111001010100;
12'd1774 : tab = 23'b00011001000100110011111;
12'd1775 : tab = 23'b00011001000010011101010;
12'd1776 : tab = 23'b00011001000000000110110;
12'd1777 : tab = 23'b00011000111101110000011;
12'd1778 : tab = 23'b00011000111011011010000;
12'd1779 : tab = 23'b00011000111001000011101;
12'd1780 : tab = 23'b00011000110110101101010;
12'd1781 : tab = 23'b00011000110100010111001;
12'd1782 : tab = 23'b00011000110010000001000;
12'd1783 : tab = 23'b00011000101111101011000;
12'd1784 : tab = 23'b00011000101101010100111;
12'd1785 : tab = 23'b00011000101010111111000;
12'd1786 : tab = 23'b00011000101000101001000;
12'd1787 : tab = 23'b00011000100110010011001;
12'd1788 : tab = 23'b00011000100011111101010;
12'd1789 : tab = 23'b00011000100001100111100;
12'd1790 : tab = 23'b00011000011111010001111;
12'd1791 : tab = 23'b00011000011100111100010;
12'd1792 : tab = 23'b00011000011010100110101;
12'd1793 : tab = 23'b00011000011000010001010;
12'd1794 : tab = 23'b00011000010101111011110;
12'd1795 : tab = 23'b00011000010011100110010;
12'd1796 : tab = 23'b00011000010001010001000;
12'd1797 : tab = 23'b00011000001110111011110;
12'd1798 : tab = 23'b00011000001100100110100;
12'd1799 : tab = 23'b00011000001010010001011;
12'd1800 : tab = 23'b00011000000111111100010;
12'd1801 : tab = 23'b00011000000101100111010;
12'd1802 : tab = 23'b00011000000011010010010;
12'd1803 : tab = 23'b00011000000000111101011;
12'd1804 : tab = 23'b00010111111110101000100;
12'd1805 : tab = 23'b00010111111100010011110;
12'd1806 : tab = 23'b00010111111001111110111;
12'd1807 : tab = 23'b00010111110111101010010;
12'd1808 : tab = 23'b00010111110101010101101;
12'd1809 : tab = 23'b00010111110011000001000;
12'd1810 : tab = 23'b00010111110000101100100;
12'd1811 : tab = 23'b00010111101110011000000;
12'd1812 : tab = 23'b00010111101100000011101;
12'd1813 : tab = 23'b00010111101001101111010;
12'd1814 : tab = 23'b00010111100111011011000;
12'd1815 : tab = 23'b00010111100101000110110;
12'd1816 : tab = 23'b00010111100010110010100;
12'd1817 : tab = 23'b00010111100000011110100;
12'd1818 : tab = 23'b00010111011110001010011;
12'd1819 : tab = 23'b00010111011011110110100;
12'd1820 : tab = 23'b00010111011001100010100;
12'd1821 : tab = 23'b00010111010111001110101;
12'd1822 : tab = 23'b00010111010100111010110;
12'd1823 : tab = 23'b00010111010010100111000;
12'd1824 : tab = 23'b00010111010000010011010;
12'd1825 : tab = 23'b00010111001101111111110;
12'd1826 : tab = 23'b00010111001011101100000;
12'd1827 : tab = 23'b00010111001001011000100;
12'd1828 : tab = 23'b00010111000111000101000;
12'd1829 : tab = 23'b00010111000100110001100;
12'd1830 : tab = 23'b00010111000010011110010;
12'd1831 : tab = 23'b00010111000000001010111;
12'd1832 : tab = 23'b00010110111101110111110;
12'd1833 : tab = 23'b00010110111011100100011;
12'd1834 : tab = 23'b00010110111001010001010;
12'd1835 : tab = 23'b00010110110110111110010;
12'd1836 : tab = 23'b00010110110100101011001;
12'd1837 : tab = 23'b00010110110010011000001;
12'd1838 : tab = 23'b00010110110000000101010;
12'd1839 : tab = 23'b00010110101101110010011;
12'd1840 : tab = 23'b00010110101011011111100;
12'd1841 : tab = 23'b00010110101001001100111;
12'd1842 : tab = 23'b00010110100110111010001;
12'd1843 : tab = 23'b00010110100100100111101;
12'd1844 : tab = 23'b00010110100010010100111;
12'd1845 : tab = 23'b00010110100000000010100;
12'd1846 : tab = 23'b00010110011101110000000;
12'd1847 : tab = 23'b00010110011011011101100;
12'd1848 : tab = 23'b00010110011001001011001;
12'd1849 : tab = 23'b00010110010110111000111;
12'd1850 : tab = 23'b00010110010100100110101;
12'd1851 : tab = 23'b00010110010010010100100;
12'd1852 : tab = 23'b00010110010000000010011;
12'd1853 : tab = 23'b00010110001101110000010;
12'd1854 : tab = 23'b00010110001011011110010;
12'd1855 : tab = 23'b00010110001001001100011;
12'd1856 : tab = 23'b00010110000110111010100;
12'd1857 : tab = 23'b00010110000100101000101;
12'd1858 : tab = 23'b00010110000010010110110;
12'd1859 : tab = 23'b00010110000000000101000;
12'd1860 : tab = 23'b00010101111101110011100;
12'd1861 : tab = 23'b00010101111011100001110;
12'd1862 : tab = 23'b00010101111001010000001;
12'd1863 : tab = 23'b00010101110110111110101;
12'd1864 : tab = 23'b00010101110100101101010;
12'd1865 : tab = 23'b00010101110010011011110;
12'd1866 : tab = 23'b00010101110000001010100;
12'd1867 : tab = 23'b00010101101101111001001;
12'd1868 : tab = 23'b00010101101011101000000;
12'd1869 : tab = 23'b00010101101001010110110;
12'd1870 : tab = 23'b00010101100111000101100;
12'd1871 : tab = 23'b00010101100100110100101;
12'd1872 : tab = 23'b00010101100010100011100;
12'd1873 : tab = 23'b00010101100000010010100;
12'd1874 : tab = 23'b00010101011110000001110;
12'd1875 : tab = 23'b00010101011011110000111;
12'd1876 : tab = 23'b00010101011001100000001;
12'd1877 : tab = 23'b00010101010111001111011;
12'd1878 : tab = 23'b00010101010100111110101;
12'd1879 : tab = 23'b00010101010010101110000;
12'd1880 : tab = 23'b00010101010000011101100;
12'd1881 : tab = 23'b00010101001110001101000;
12'd1882 : tab = 23'b00010101001011111100100;
12'd1883 : tab = 23'b00010101001001101100010;
12'd1884 : tab = 23'b00010101000111011011110;
12'd1885 : tab = 23'b00010101000101001011100;
12'd1886 : tab = 23'b00010101000010111011010;
12'd1887 : tab = 23'b00010101000000101011000;
12'd1888 : tab = 23'b00010100111110011011000;
12'd1889 : tab = 23'b00010100111100001010111;
12'd1890 : tab = 23'b00010100111001111010111;
12'd1891 : tab = 23'b00010100110111101010111;
12'd1892 : tab = 23'b00010100110101011011000;
12'd1893 : tab = 23'b00010100110011001011000;
12'd1894 : tab = 23'b00010100110000111011010;
12'd1895 : tab = 23'b00010100101110101011101;
12'd1896 : tab = 23'b00010100101100011011111;
12'd1897 : tab = 23'b00010100101010001100010;
12'd1898 : tab = 23'b00010100100111111100110;
12'd1899 : tab = 23'b00010100100101101101001;
12'd1900 : tab = 23'b00010100100011011101110;
12'd1901 : tab = 23'b00010100100001001110010;
12'd1902 : tab = 23'b00010100011110111111000;
12'd1903 : tab = 23'b00010100011100101111100;
12'd1904 : tab = 23'b00010100011010100000010;
12'd1905 : tab = 23'b00010100011000010001010;
12'd1906 : tab = 23'b00010100010110000010000;
12'd1907 : tab = 23'b00010100010011110011000;
12'd1908 : tab = 23'b00010100010001100011111;
12'd1909 : tab = 23'b00010100001111010101000;
12'd1910 : tab = 23'b00010100001101000110000;
12'd1911 : tab = 23'b00010100001010110111000;
12'd1912 : tab = 23'b00010100001000101000010;
12'd1913 : tab = 23'b00010100000110011001100;
12'd1914 : tab = 23'b00010100000100001010110;
12'd1915 : tab = 23'b00010100000001111100001;
12'd1916 : tab = 23'b00010011111111101101101;
12'd1917 : tab = 23'b00010011111101011111000;
12'd1918 : tab = 23'b00010011111011010000101;
12'd1919 : tab = 23'b00010011111001000010001;
12'd1920 : tab = 23'b00010011110110110011110;
12'd1921 : tab = 23'b00010011110100100101011;
12'd1922 : tab = 23'b00010011110010010111001;
12'd1923 : tab = 23'b00010011110000001000111;
12'd1924 : tab = 23'b00010011101101111010110;
12'd1925 : tab = 23'b00010011101011101100101;
12'd1926 : tab = 23'b00010011101001011110100;
12'd1927 : tab = 23'b00010011100111010000100;
12'd1928 : tab = 23'b00010011100101000010101;
12'd1929 : tab = 23'b00010011100010110100101;
12'd1930 : tab = 23'b00010011100000100110110;
12'd1931 : tab = 23'b00010011011110011001000;
12'd1932 : tab = 23'b00010011011100001011010;
12'd1933 : tab = 23'b00010011011001111101100;
12'd1934 : tab = 23'b00010011010111110000000;
12'd1935 : tab = 23'b00010011010101100010011;
12'd1936 : tab = 23'b00010011010011010100110;
12'd1937 : tab = 23'b00010011010001000111010;
12'd1938 : tab = 23'b00010011001110111001111;
12'd1939 : tab = 23'b00010011001100101100100;
12'd1940 : tab = 23'b00010011001010011111010;
12'd1941 : tab = 23'b00010011001000010010000;
12'd1942 : tab = 23'b00010011000110000100110;
12'd1943 : tab = 23'b00010011000011110111100;
12'd1944 : tab = 23'b00010011000001101010100;
12'd1945 : tab = 23'b00010010111111011101011;
12'd1946 : tab = 23'b00010010111101010000011;
12'd1947 : tab = 23'b00010010111011000011011;
12'd1948 : tab = 23'b00010010111000110110100;
12'd1949 : tab = 23'b00010010110110101001110;
12'd1950 : tab = 23'b00010010110100011101000;
12'd1951 : tab = 23'b00010010110010010000010;
12'd1952 : tab = 23'b00010010110000000011101;
12'd1953 : tab = 23'b00010010101101110111000;
12'd1954 : tab = 23'b00010010101011101010011;
12'd1955 : tab = 23'b00010010101001011101110;
12'd1956 : tab = 23'b00010010100111010001011;
12'd1957 : tab = 23'b00010010100101000101000;
12'd1958 : tab = 23'b00010010100010111000101;
12'd1959 : tab = 23'b00010010100000101100010;
12'd1960 : tab = 23'b00010010011110100000000;
12'd1961 : tab = 23'b00010010011100010011110;
12'd1962 : tab = 23'b00010010011010000111110;
12'd1963 : tab = 23'b00010010010111111011100;
12'd1964 : tab = 23'b00010010010101101111100;
12'd1965 : tab = 23'b00010010010011100011100;
12'd1966 : tab = 23'b00010010010001010111100;
12'd1967 : tab = 23'b00010010001111001011101;
12'd1968 : tab = 23'b00010010001100111111110;
12'd1969 : tab = 23'b00010010001010110100000;
12'd1970 : tab = 23'b00010010001000101000010;
12'd1971 : tab = 23'b00010010000110011100101;
12'd1972 : tab = 23'b00010010000100010001000;
12'd1973 : tab = 23'b00010010000010000101011;
12'd1974 : tab = 23'b00010001111111111010000;
12'd1975 : tab = 23'b00010001111101101110100;
12'd1976 : tab = 23'b00010001111011100011000;
12'd1977 : tab = 23'b00010001111001010111101;
12'd1978 : tab = 23'b00010001110111001100010;
12'd1979 : tab = 23'b00010001110101000001000;
12'd1980 : tab = 23'b00010001110010110101110;
12'd1981 : tab = 23'b00010001110000101010100;
12'd1982 : tab = 23'b00010001101110011111100;
12'd1983 : tab = 23'b00010001101100010100011;
12'd1984 : tab = 23'b00010001101010001001011;
12'd1985 : tab = 23'b00010001100111111110100;
12'd1986 : tab = 23'b00010001100101110011100;
12'd1987 : tab = 23'b00010001100011101000110;
12'd1988 : tab = 23'b00010001100001011101111;
12'd1989 : tab = 23'b00010001011111010011010;
12'd1990 : tab = 23'b00010001011101001000100;
12'd1991 : tab = 23'b00010001011010111101110;
12'd1992 : tab = 23'b00010001011000110011010;
12'd1993 : tab = 23'b00010001010110101000101;
12'd1994 : tab = 23'b00010001010100011110001;
12'd1995 : tab = 23'b00010001010010010011110;
12'd1996 : tab = 23'b00010001010000001001010;
12'd1997 : tab = 23'b00010001001101111111000;
12'd1998 : tab = 23'b00010001001011110100110;
12'd1999 : tab = 23'b00010001001001101010100;
12'd2000 : tab = 23'b00010001000111100000010;
12'd2001 : tab = 23'b00010001000101010110001;
12'd2002 : tab = 23'b00010001000011001100000;
12'd2003 : tab = 23'b00010001000001000010000;
12'd2004 : tab = 23'b00010000111110111000000;
12'd2005 : tab = 23'b00010000111100101110001;
12'd2006 : tab = 23'b00010000111010100100010;
12'd2007 : tab = 23'b00010000111000011010011;
12'd2008 : tab = 23'b00010000110110010000100;
12'd2009 : tab = 23'b00010000110100000111000;
12'd2010 : tab = 23'b00010000110001111101010;
12'd2011 : tab = 23'b00010000101111110011110;
12'd2012 : tab = 23'b00010000101101101010000;
12'd2013 : tab = 23'b00010000101011100000100;
12'd2014 : tab = 23'b00010000101001010111000;
12'd2015 : tab = 23'b00010000100111001101100;
12'd2016 : tab = 23'b00010000100101000100010;
12'd2017 : tab = 23'b00010000100010111011000;
12'd2018 : tab = 23'b00010000100000110001101;
12'd2019 : tab = 23'b00010000011110101000011;
12'd2020 : tab = 23'b00010000011100011111010;
12'd2021 : tab = 23'b00010000011010010110001;
12'd2022 : tab = 23'b00010000011000001101001;
12'd2023 : tab = 23'b00010000010110000100001;
12'd2024 : tab = 23'b00010000010011111011000;
12'd2025 : tab = 23'b00010000010001110010001;
12'd2026 : tab = 23'b00010000001111101001010;
12'd2027 : tab = 23'b00010000001101100000100;
12'd2028 : tab = 23'b00010000001011010111110;
12'd2029 : tab = 23'b00010000001001001111000;
12'd2030 : tab = 23'b00010000000111000110011;
12'd2031 : tab = 23'b00010000000100111101110;
12'd2032 : tab = 23'b00010000000010110101010;
12'd2033 : tab = 23'b00010000000000101100110;
12'd2034 : tab = 23'b00001111111110100100010;
12'd2035 : tab = 23'b00001111111100011011110;
12'd2036 : tab = 23'b00001111111010010011011;
12'd2037 : tab = 23'b00001111111000001011000;
12'd2038 : tab = 23'b00001111110110000010111;
12'd2039 : tab = 23'b00001111110011111010101;
12'd2040 : tab = 23'b00001111110001110010100;
12'd2041 : tab = 23'b00001111101111101010011;
12'd2042 : tab = 23'b00001111101101100010010;
12'd2043 : tab = 23'b00001111101011011010010;
12'd2044 : tab = 23'b00001111101001010010010;
12'd2045 : tab = 23'b00001111100111001010100;
12'd2046 : tab = 23'b00001111100101000010100;
12'd2047 : tab = 23'b00001111100010111010110;
12'd2048 : tab = 23'b00001111011111101111001;
12'd2049 : tab = 23'b00001111011011011111110;
12'd2050 : tab = 23'b00001111010111010000110;
12'd2051 : tab = 23'b00001111010011000001110;
12'd2052 : tab = 23'b00001111001110110011000;
12'd2053 : tab = 23'b00001111001010100100100;
12'd2054 : tab = 23'b00001111000110010110001;
12'd2055 : tab = 23'b00001111000010001000000;
12'd2056 : tab = 23'b00001110111101111010000;
12'd2057 : tab = 23'b00001110111001101100010;
12'd2058 : tab = 23'b00001110110101011110110;
12'd2059 : tab = 23'b00001110110001010001011;
12'd2060 : tab = 23'b00001110101101000100010;
12'd2061 : tab = 23'b00001110101000110111010;
12'd2062 : tab = 23'b00001110100100101010100;
12'd2063 : tab = 23'b00001110100000011101111;
12'd2064 : tab = 23'b00001110011100010001100;
12'd2065 : tab = 23'b00001110011000000101011;
12'd2066 : tab = 23'b00001110010011111001010;
12'd2067 : tab = 23'b00001110001111101101100;
12'd2068 : tab = 23'b00001110001011100010000;
12'd2069 : tab = 23'b00001110000111010110100;
12'd2070 : tab = 23'b00001110000011001011010;
12'd2071 : tab = 23'b00001101111111000000011;
12'd2072 : tab = 23'b00001101111010110101100;
12'd2073 : tab = 23'b00001101110110101010110;
12'd2074 : tab = 23'b00001101110010100000011;
12'd2075 : tab = 23'b00001101101110010110001;
12'd2076 : tab = 23'b00001101101010001100000;
12'd2077 : tab = 23'b00001101100110000010010;
12'd2078 : tab = 23'b00001101100001111000101;
12'd2079 : tab = 23'b00001101011101101111001;
12'd2080 : tab = 23'b00001101011001100101110;
12'd2081 : tab = 23'b00001101010101011100110;
12'd2082 : tab = 23'b00001101010001010011110;
12'd2083 : tab = 23'b00001101001101001011000;
12'd2084 : tab = 23'b00001101001001000010101;
12'd2085 : tab = 23'b00001101000100111010010;
12'd2086 : tab = 23'b00001101000000110010001;
12'd2087 : tab = 23'b00001100111100101010001;
12'd2088 : tab = 23'b00001100111000100010011;
12'd2089 : tab = 23'b00001100110100011010111;
12'd2090 : tab = 23'b00001100110000010011100;
12'd2091 : tab = 23'b00001100101100001100010;
12'd2092 : tab = 23'b00001100101000000101010;
12'd2093 : tab = 23'b00001100100011111110100;
12'd2094 : tab = 23'b00001100011111110111110;
12'd2095 : tab = 23'b00001100011011110001010;
12'd2096 : tab = 23'b00001100010111101011000;
12'd2097 : tab = 23'b00001100010011100101000;
12'd2098 : tab = 23'b00001100001111011111001;
12'd2099 : tab = 23'b00001100001011011001011;
12'd2100 : tab = 23'b00001100000111010100000;
12'd2101 : tab = 23'b00001100000011001110100;
12'd2102 : tab = 23'b00001011111111001001100;
12'd2103 : tab = 23'b00001011111011000100100;
12'd2104 : tab = 23'b00001011110110111111110;
12'd2105 : tab = 23'b00001011110010111011001;
12'd2106 : tab = 23'b00001011101110110110111;
12'd2107 : tab = 23'b00001011101010110010101;
12'd2108 : tab = 23'b00001011100110101110100;
12'd2109 : tab = 23'b00001011100010101010110;
12'd2110 : tab = 23'b00001011011110100111001;
12'd2111 : tab = 23'b00001011011010100011110;
12'd2112 : tab = 23'b00001011010110100000011;
12'd2113 : tab = 23'b00001011010010011101010;
12'd2114 : tab = 23'b00001011001110011010010;
12'd2115 : tab = 23'b00001011001010010111101;
12'd2116 : tab = 23'b00001011000110010101001;
12'd2117 : tab = 23'b00001011000010010010101;
12'd2118 : tab = 23'b00001010111110010000100;
12'd2119 : tab = 23'b00001010111010001110100;
12'd2120 : tab = 23'b00001010110110001100110;
12'd2121 : tab = 23'b00001010110010001011000;
12'd2122 : tab = 23'b00001010101110001001100;
12'd2123 : tab = 23'b00001010101010001000010;
12'd2124 : tab = 23'b00001010100110000111010;
12'd2125 : tab = 23'b00001010100010000110011;
12'd2126 : tab = 23'b00001010011110000101110;
12'd2127 : tab = 23'b00001010011010000101000;
12'd2128 : tab = 23'b00001010010110000100110;
12'd2129 : tab = 23'b00001010010010000100100;
12'd2130 : tab = 23'b00001010001110000100100;
12'd2131 : tab = 23'b00001010001010000100110;
12'd2132 : tab = 23'b00001010000110000101001;
12'd2133 : tab = 23'b00001010000010000101100;
12'd2134 : tab = 23'b00001001111110000110011;
12'd2135 : tab = 23'b00001001111010000111010;
12'd2136 : tab = 23'b00001001110110001000011;
12'd2137 : tab = 23'b00001001110010001001100;
12'd2138 : tab = 23'b00001001101110001011000;
12'd2139 : tab = 23'b00001001101010001100101;
12'd2140 : tab = 23'b00001001100110001110100;
12'd2141 : tab = 23'b00001001100010010000011;
12'd2142 : tab = 23'b00001001011110010010100;
12'd2143 : tab = 23'b00001001011010010100110;
12'd2144 : tab = 23'b00001001010110010111011;
12'd2145 : tab = 23'b00001001010010011010000;
12'd2146 : tab = 23'b00001001001110011100111;
12'd2147 : tab = 23'b00001001001010100000000;
12'd2148 : tab = 23'b00001001000110100011010;
12'd2149 : tab = 23'b00001001000010100110100;
12'd2150 : tab = 23'b00001000111110101010000;
12'd2151 : tab = 23'b00001000111010101101111;
12'd2152 : tab = 23'b00001000110110110001110;
12'd2153 : tab = 23'b00001000110010110101111;
12'd2154 : tab = 23'b00001000101110111010000;
12'd2155 : tab = 23'b00001000101010111110101;
12'd2156 : tab = 23'b00001000100111000011010;
12'd2157 : tab = 23'b00001000100011001000000;
12'd2158 : tab = 23'b00001000011111001100111;
12'd2159 : tab = 23'b00001000011011010010000;
12'd2160 : tab = 23'b00001000010111010111011;
12'd2161 : tab = 23'b00001000010011011100110;
12'd2162 : tab = 23'b00001000001111100010100;
12'd2163 : tab = 23'b00001000001011101000011;
12'd2164 : tab = 23'b00001000000111101110011;
12'd2165 : tab = 23'b00001000000011110100100;
12'd2166 : tab = 23'b00000111111111111011000;
12'd2167 : tab = 23'b00000111111100000001011;
12'd2168 : tab = 23'b00000111111000001000010;
12'd2169 : tab = 23'b00000111110100001111000;
12'd2170 : tab = 23'b00000111110000010110000;
12'd2171 : tab = 23'b00000111101100011101010;
12'd2172 : tab = 23'b00000111101000100100101;
12'd2173 : tab = 23'b00000111100100101100001;
12'd2174 : tab = 23'b00000111100000110011111;
12'd2175 : tab = 23'b00000111011100111011110;
12'd2176 : tab = 23'b00000111011001000100000;
12'd2177 : tab = 23'b00000111010101001100010;
12'd2178 : tab = 23'b00000111010001010100100;
12'd2179 : tab = 23'b00000111001101011101001;
12'd2180 : tab = 23'b00000111001001100110000;
12'd2181 : tab = 23'b00000111000101101110110;
12'd2182 : tab = 23'b00000111000001110111111;
12'd2183 : tab = 23'b00000110111110000001001;
12'd2184 : tab = 23'b00000110111010001010101;
12'd2185 : tab = 23'b00000110110110010100010;
12'd2186 : tab = 23'b00000110110010011110000;
12'd2187 : tab = 23'b00000110101110101000000;
12'd2188 : tab = 23'b00000110101010110010000;
12'd2189 : tab = 23'b00000110100110111100011;
12'd2190 : tab = 23'b00000110100011000110110;
12'd2191 : tab = 23'b00000110011111010001010;
12'd2192 : tab = 23'b00000110011011011100010;
12'd2193 : tab = 23'b00000110010111100111001;
12'd2194 : tab = 23'b00000110010011110010010;
12'd2195 : tab = 23'b00000110001111111101101;
12'd2196 : tab = 23'b00000110001100001001000;
12'd2197 : tab = 23'b00000110001000010100101;
12'd2198 : tab = 23'b00000110000100100000011;
12'd2199 : tab = 23'b00000110000000101100011;
12'd2200 : tab = 23'b00000101111100111000100;
12'd2201 : tab = 23'b00000101111001000100110;
12'd2202 : tab = 23'b00000101110101010001010;
12'd2203 : tab = 23'b00000101110001011101110;
12'd2204 : tab = 23'b00000101101101101010100;
12'd2205 : tab = 23'b00000101101001110111100;
12'd2206 : tab = 23'b00000101100110000100101;
12'd2207 : tab = 23'b00000101100010010010000;
12'd2208 : tab = 23'b00000101011110011111011;
12'd2209 : tab = 23'b00000101011010101101000;
12'd2210 : tab = 23'b00000101010110111010110;
12'd2211 : tab = 23'b00000101010011001000110;
12'd2212 : tab = 23'b00000101001111010110111;
12'd2213 : tab = 23'b00000101001011100101001;
12'd2214 : tab = 23'b00000101000111110011100;
12'd2215 : tab = 23'b00000101000100000010010;
12'd2216 : tab = 23'b00000101000000010000111;
12'd2217 : tab = 23'b00000100111100011111110;
12'd2218 : tab = 23'b00000100111000101110111;
12'd2219 : tab = 23'b00000100110100111110000;
12'd2220 : tab = 23'b00000100110001001101100;
12'd2221 : tab = 23'b00000100101101011101001;
12'd2222 : tab = 23'b00000100101001101100110;
12'd2223 : tab = 23'b00000100100101111100110;
12'd2224 : tab = 23'b00000100100010001100110;
12'd2225 : tab = 23'b00000100011110011101000;
12'd2226 : tab = 23'b00000100011010101101011;
12'd2227 : tab = 23'b00000100010110111101111;
12'd2228 : tab = 23'b00000100010011001110101;
12'd2229 : tab = 23'b00000100001111011111011;
12'd2230 : tab = 23'b00000100001011110000100;
12'd2231 : tab = 23'b00000100001000000001101;
12'd2232 : tab = 23'b00000100000100010011000;
12'd2233 : tab = 23'b00000100000000100100100;
12'd2234 : tab = 23'b00000011111100110110001;
12'd2235 : tab = 23'b00000011111001001000000;
12'd2236 : tab = 23'b00000011110101011010000;
12'd2237 : tab = 23'b00000011110001101100001;
12'd2238 : tab = 23'b00000011101101111110011;
12'd2239 : tab = 23'b00000011101010010000111;
12'd2240 : tab = 23'b00000011100110100011100;
12'd2241 : tab = 23'b00000011100010110110011;
12'd2242 : tab = 23'b00000011011111001001010;
12'd2243 : tab = 23'b00000011011011011100011;
12'd2244 : tab = 23'b00000011010111101111101;
12'd2245 : tab = 23'b00000011010100000011000;
12'd2246 : tab = 23'b00000011010000010110100;
12'd2247 : tab = 23'b00000011001100101010010;
12'd2248 : tab = 23'b00000011001000111110010;
12'd2249 : tab = 23'b00000011000101010010010;
12'd2250 : tab = 23'b00000011000001100110100;
12'd2251 : tab = 23'b00000010111101111010110;
12'd2252 : tab = 23'b00000010111010001111010;
12'd2253 : tab = 23'b00000010110110100100000;
12'd2254 : tab = 23'b00000010110010111000111;
12'd2255 : tab = 23'b00000010101111001110000;
12'd2256 : tab = 23'b00000010101011100011000;
12'd2257 : tab = 23'b00000010100111111000011;
12'd2258 : tab = 23'b00000010100100001101110;
12'd2259 : tab = 23'b00000010100000100011010;
12'd2260 : tab = 23'b00000010011100111001001;
12'd2261 : tab = 23'b00000010011001001111000;
12'd2262 : tab = 23'b00000010010101100101001;
12'd2263 : tab = 23'b00000010010001111011011;
12'd2264 : tab = 23'b00000010001110010001110;
12'd2265 : tab = 23'b00000010001010101000010;
12'd2266 : tab = 23'b00000010000110111111000;
12'd2267 : tab = 23'b00000010000011010101111;
12'd2268 : tab = 23'b00000001111111101100111;
12'd2269 : tab = 23'b00000001111100000100000;
12'd2270 : tab = 23'b00000001111000011011010;
12'd2271 : tab = 23'b00000001110100110010110;
12'd2272 : tab = 23'b00000001110001001010011;
12'd2273 : tab = 23'b00000001101101100010010;
12'd2274 : tab = 23'b00000001101001111010000;
12'd2275 : tab = 23'b00000001100110010010001;
12'd2276 : tab = 23'b00000001100010101010011;
12'd2277 : tab = 23'b00000001011111000010110;
12'd2278 : tab = 23'b00000001011011011011100;
12'd2279 : tab = 23'b00000001010111110100000;
12'd2280 : tab = 23'b00000001010100001100111;
12'd2281 : tab = 23'b00000001010000100101111;
12'd2282 : tab = 23'b00000001001100111111000;
12'd2283 : tab = 23'b00000001001001011000010;
12'd2284 : tab = 23'b00000001000101110001110;
12'd2285 : tab = 23'b00000001000010001011011;
12'd2286 : tab = 23'b00000000111110100101001;
12'd2287 : tab = 23'b00000000111010111111000;
12'd2288 : tab = 23'b00000000110111011001000;
12'd2289 : tab = 23'b00000000110011110011010;
12'd2290 : tab = 23'b00000000110000001101101;
12'd2291 : tab = 23'b00000000101100101000001;
12'd2292 : tab = 23'b00000000101001000010110;
12'd2293 : tab = 23'b00000000100101011101100;
12'd2294 : tab = 23'b00000000100001111000100;
12'd2295 : tab = 23'b00000000011110010011101;
12'd2296 : tab = 23'b00000000011010101110111;
12'd2297 : tab = 23'b00000000010111001010010;
12'd2298 : tab = 23'b00000000010011100101111;
12'd2299 : tab = 23'b00000000010000000001100;
12'd2300 : tab = 23'b00000000001100011101011;
12'd2301 : tab = 23'b00000000001000111001011;
12'd2302 : tab = 23'b00000000000101010101100;
12'd2303 : tab = 23'b00000000000001110010000;
12'd2304 : tab = 23'b11111111111100011100101;
12'd2305 : tab = 23'b11111111110101010101110;
12'd2306 : tab = 23'b11111111101110001111010;
12'd2307 : tab = 23'b11111111100111001001001;
12'd2308 : tab = 23'b11111111100000000011000;
12'd2309 : tab = 23'b11111111011000111101100;
12'd2310 : tab = 23'b11111111010001111000010;
12'd2311 : tab = 23'b11111111001010110011000;
12'd2312 : tab = 23'b11111111000011101110010;
12'd2313 : tab = 23'b11111110111100101010000;
12'd2314 : tab = 23'b11111110110101100101110;
12'd2315 : tab = 23'b11111110101110100001111;
12'd2316 : tab = 23'b11111110100111011110011;
12'd2317 : tab = 23'b11111110100000011010111;
12'd2318 : tab = 23'b11111110011001011000001;
12'd2319 : tab = 23'b11111110010010010101011;
12'd2320 : tab = 23'b11111110001011010011000;
12'd2321 : tab = 23'b11111110000100010000101;
12'd2322 : tab = 23'b11111101111101001111000;
12'd2323 : tab = 23'b11111101110110001101011;
12'd2324 : tab = 23'b11111101101111001100001;
12'd2325 : tab = 23'b11111101101000001011010;
12'd2326 : tab = 23'b11111101100001001010011;
12'd2327 : tab = 23'b11111101011010001010010;
12'd2328 : tab = 23'b11111101010011001010001;
12'd2329 : tab = 23'b11111101001100001010011;
12'd2330 : tab = 23'b11111101000101001010101;
12'd2331 : tab = 23'b11111100111110001011100;
12'd2332 : tab = 23'b11111100110111001100100;
12'd2333 : tab = 23'b11111100110000001101110;
12'd2334 : tab = 23'b11111100101001001111011;
12'd2335 : tab = 23'b11111100100010010001100;
12'd2336 : tab = 23'b11111100011011010011101;
12'd2337 : tab = 23'b11111100010100010110001;
12'd2338 : tab = 23'b11111100001101011001000;
12'd2339 : tab = 23'b11111100000110011011111;
12'd2340 : tab = 23'b11111011111111011111010;
12'd2341 : tab = 23'b11111011111000100011001;
12'd2342 : tab = 23'b11111011110001100111000;
12'd2343 : tab = 23'b11111011101010101011001;
12'd2344 : tab = 23'b11111011100011101111100;
12'd2345 : tab = 23'b11111011011100110100100;
12'd2346 : tab = 23'b11111011010101111001011;
12'd2347 : tab = 23'b11111011001110111110111;
12'd2348 : tab = 23'b11111011001000000100011;
12'd2349 : tab = 23'b11111011000001001010010;
12'd2350 : tab = 23'b11111010111010010000100;
12'd2351 : tab = 23'b11111010110011010111000;
12'd2352 : tab = 23'b11111010101100011101110;
12'd2353 : tab = 23'b11111010100101100100110;
12'd2354 : tab = 23'b11111010011110101100001;
12'd2355 : tab = 23'b11111010010111110011100;
12'd2356 : tab = 23'b11111010010000111011101;
12'd2357 : tab = 23'b11111010001010000011110;
12'd2358 : tab = 23'b11111010000011001100010;
12'd2359 : tab = 23'b11111001111100010100110;
12'd2360 : tab = 23'b11111001110101011101110;
12'd2361 : tab = 23'b11111001101110100110111;
12'd2362 : tab = 23'b11111001100111110000100;
12'd2363 : tab = 23'b11111001100000111010100;
12'd2364 : tab = 23'b11111001011010000100100;
12'd2365 : tab = 23'b11111001010011001110111;
12'd2366 : tab = 23'b11111001001100011001101;
12'd2367 : tab = 23'b11111001000101100100011;
12'd2368 : tab = 23'b11111000111110101111110;
12'd2369 : tab = 23'b11111000110111111011010;
12'd2370 : tab = 23'b11111000110001000111000;
12'd2371 : tab = 23'b11111000101010010011001;
12'd2372 : tab = 23'b11111000100011011111011;
12'd2373 : tab = 23'b11111000011100101100000;
12'd2374 : tab = 23'b11111000010101111000110;
12'd2375 : tab = 23'b11111000001111000110000;
12'd2376 : tab = 23'b11111000001000010011011;
12'd2377 : tab = 23'b11111000000001100001001;
12'd2378 : tab = 23'b11110111111010101111000;
12'd2379 : tab = 23'b11110111110011111101011;
12'd2380 : tab = 23'b11110111101101001011111;
12'd2381 : tab = 23'b11110111100110011010100;
12'd2382 : tab = 23'b11110111011111101001101;
12'd2383 : tab = 23'b11110111011000111000111;
12'd2384 : tab = 23'b11110111010010001000100;
12'd2385 : tab = 23'b11110111001011011000100;
12'd2386 : tab = 23'b11110111000100101000100;
12'd2387 : tab = 23'b11110110111101111000111;
12'd2388 : tab = 23'b11110110110111001001101;
12'd2389 : tab = 23'b11110110110000011010110;
12'd2390 : tab = 23'b11110110101001101011111;
12'd2391 : tab = 23'b11110110100010111101011;
12'd2392 : tab = 23'b11110110011100001111010;
12'd2393 : tab = 23'b11110110010101100001001;
12'd2394 : tab = 23'b11110110001110110011011;
12'd2395 : tab = 23'b11110110001000000110000;
12'd2396 : tab = 23'b11110110000001011001000;
12'd2397 : tab = 23'b11110101111010101100000;
12'd2398 : tab = 23'b11110101110011111111011;
12'd2399 : tab = 23'b11110101101101010011001;
12'd2400 : tab = 23'b11110101100110100110111;
12'd2401 : tab = 23'b11110101011111111011010;
12'd2402 : tab = 23'b11110101011001001111100;
12'd2403 : tab = 23'b11110101010010100100011;
12'd2404 : tab = 23'b11110101001011111001010;
12'd2405 : tab = 23'b11110101000101001110100;
12'd2406 : tab = 23'b11110100111110100100001;
12'd2407 : tab = 23'b11110100110111111010000;
12'd2408 : tab = 23'b11110100110001010000000;
12'd2409 : tab = 23'b11110100101010100110010;
12'd2410 : tab = 23'b11110100100011111100111;
12'd2411 : tab = 23'b11110100011101010011101;
12'd2412 : tab = 23'b11110100010110101010110;
12'd2413 : tab = 23'b11110100010000000010010;
12'd2414 : tab = 23'b11110100001001011010000;
12'd2415 : tab = 23'b11110100000010110001101;
12'd2416 : tab = 23'b11110011111100001001111;
12'd2417 : tab = 23'b11110011110101100010010;
12'd2418 : tab = 23'b11110011101110111011001;
12'd2419 : tab = 23'b11110011101000010100001;
12'd2420 : tab = 23'b11110011100001101101001;
12'd2421 : tab = 23'b11110011011011000110110;
12'd2422 : tab = 23'b11110011010100100000100;
12'd2423 : tab = 23'b11110011001101111010011;
12'd2424 : tab = 23'b11110011000111010100110;
12'd2425 : tab = 23'b11110011000000101111000;
12'd2426 : tab = 23'b11110010111010001001111;
12'd2427 : tab = 23'b11110010110011100101001;
12'd2428 : tab = 23'b11110010101101000000011;
12'd2429 : tab = 23'b11110010100110011100000;
12'd2430 : tab = 23'b11110010011111110111110;
12'd2431 : tab = 23'b11110010011001010011101;
12'd2432 : tab = 23'b11110010010010110000000;
12'd2433 : tab = 23'b11110010001100001100110;
12'd2434 : tab = 23'b11110010000101101001100;
12'd2435 : tab = 23'b11110001111111000110110;
12'd2436 : tab = 23'b11110001111000100100001;
12'd2437 : tab = 23'b11110001110010000001101;
12'd2438 : tab = 23'b11110001101011011111100;
12'd2439 : tab = 23'b11110001100100111101110;
12'd2440 : tab = 23'b11110001011110011100010;
12'd2441 : tab = 23'b11110001010111111010110;
12'd2442 : tab = 23'b11110001010001011001110;
12'd2443 : tab = 23'b11110001001010111001000;
12'd2444 : tab = 23'b11110001000100011000011;
12'd2445 : tab = 23'b11110000111101111000001;
12'd2446 : tab = 23'b11110000110111010111111;
12'd2447 : tab = 23'b11110000110000111000010;
12'd2448 : tab = 23'b11110000101010011000100;
12'd2449 : tab = 23'b11110000100011111001011;
12'd2450 : tab = 23'b11110000011101011010010;
12'd2451 : tab = 23'b11110000010110111011100;
12'd2452 : tab = 23'b11110000010000011101000;
12'd2453 : tab = 23'b11110000001001111110110;
12'd2454 : tab = 23'b11110000000011100000110;
12'd2455 : tab = 23'b11101111111101000010110;
12'd2456 : tab = 23'b11101111110110100101010;
12'd2457 : tab = 23'b11101111110000001000000;
12'd2458 : tab = 23'b11101111101001101011000;
12'd2459 : tab = 23'b11101111100011001110010;
12'd2460 : tab = 23'b11101111011100110001110;
12'd2461 : tab = 23'b11101111010110010101100;
12'd2462 : tab = 23'b11101111001111111001011;
12'd2463 : tab = 23'b11101111001001011101110;
12'd2464 : tab = 23'b11101111000011000010010;
12'd2465 : tab = 23'b11101110111100100111000;
12'd2466 : tab = 23'b11101110110110001100000;
12'd2467 : tab = 23'b11101110101111110001010;
12'd2468 : tab = 23'b11101110101001010110101;
12'd2469 : tab = 23'b11101110100010111100011;
12'd2470 : tab = 23'b11101110011100100010100;
12'd2471 : tab = 23'b11101110010110001000101;
12'd2472 : tab = 23'b11101110001111101111001;
12'd2473 : tab = 23'b11101110001001010101110;
12'd2474 : tab = 23'b11101110000010111100111;
12'd2475 : tab = 23'b11101101111100100100001;
12'd2476 : tab = 23'b11101101110110001011100;
12'd2477 : tab = 23'b11101101101111110011011;
12'd2478 : tab = 23'b11101101101001011011011;
12'd2479 : tab = 23'b11101101100011000011011;
12'd2480 : tab = 23'b11101101011100101100000;
12'd2481 : tab = 23'b11101101010110010100110;
12'd2482 : tab = 23'b11101101001111111101101;
12'd2483 : tab = 23'b11101101001001100110110;
12'd2484 : tab = 23'b11101101000011010000010;
12'd2485 : tab = 23'b11101100111100111010000;
12'd2486 : tab = 23'b11101100110110100100000;
12'd2487 : tab = 23'b11101100110000001110010;
12'd2488 : tab = 23'b11101100101001111000100;
12'd2489 : tab = 23'b11101100100011100011001;
12'd2490 : tab = 23'b11101100011101001110001;
12'd2491 : tab = 23'b11101100010110111001010;
12'd2492 : tab = 23'b11101100010000100100110;
12'd2493 : tab = 23'b11101100001010010000010;
12'd2494 : tab = 23'b11101100000011111100010;
12'd2495 : tab = 23'b11101011111101101000100;
12'd2496 : tab = 23'b11101011110111010100110;
12'd2497 : tab = 23'b11101011110001000001100;
12'd2498 : tab = 23'b11101011101010101110011;
12'd2499 : tab = 23'b11101011100100011011100;
12'd2500 : tab = 23'b11101011011110001000110;
12'd2501 : tab = 23'b11101011010111110110100;
12'd2502 : tab = 23'b11101011010001100100001;
12'd2503 : tab = 23'b11101011001011010010001;
12'd2504 : tab = 23'b11101011000101000000100;
12'd2505 : tab = 23'b11101010111110101111000;
12'd2506 : tab = 23'b11101010111000011110000;
12'd2507 : tab = 23'b11101010110010001101000;
12'd2508 : tab = 23'b11101010101011111100010;
12'd2509 : tab = 23'b11101010100101101011110;
12'd2510 : tab = 23'b11101010011111011011100;
12'd2511 : tab = 23'b11101010011001001011100;
12'd2512 : tab = 23'b11101010010010111011110;
12'd2513 : tab = 23'b11101010001100101100000;
12'd2514 : tab = 23'b11101010000110011100110;
12'd2515 : tab = 23'b11101010000000001101101;
12'd2516 : tab = 23'b11101001111001111111000;
12'd2517 : tab = 23'b11101001110011110000011;
12'd2518 : tab = 23'b11101001101101100010001;
12'd2519 : tab = 23'b11101001100111010011111;
12'd2520 : tab = 23'b11101001100001000110000;
12'd2521 : tab = 23'b11101001011010111000010;
12'd2522 : tab = 23'b11101001010100101011000;
12'd2523 : tab = 23'b11101001001110011101111;
12'd2524 : tab = 23'b11101001001000010001000;
12'd2525 : tab = 23'b11101001000010000100010;
12'd2526 : tab = 23'b11101000111011110111110;
12'd2527 : tab = 23'b11101000110101101011101;
12'd2528 : tab = 23'b11101000101111011111101;
12'd2529 : tab = 23'b11101000101001010011101;
12'd2530 : tab = 23'b11101000100011001000011;
12'd2531 : tab = 23'b11101000011100111101001;
12'd2532 : tab = 23'b11101000010110110010000;
12'd2533 : tab = 23'b11101000010000100111010;
12'd2534 : tab = 23'b11101000001010011100100;
12'd2535 : tab = 23'b11101000000100010010010;
12'd2536 : tab = 23'b11100111111110001000000;
12'd2537 : tab = 23'b11100111110111111110010;
12'd2538 : tab = 23'b11100111110001110100110;
12'd2539 : tab = 23'b11100111101011101011010;
12'd2540 : tab = 23'b11100111100101100010010;
12'd2541 : tab = 23'b11100111011111011001000;
12'd2542 : tab = 23'b11100111011001010000011;
12'd2543 : tab = 23'b11100111010011000111110;
12'd2544 : tab = 23'b11100111001100111111100;
12'd2545 : tab = 23'b11100111000110110111101;
12'd2546 : tab = 23'b11100111000000101111110;
12'd2547 : tab = 23'b11100110111010101000010;
12'd2548 : tab = 23'b11100110110100100001000;
12'd2549 : tab = 23'b11100110101110011010000;
12'd2550 : tab = 23'b11100110101000010010111;
12'd2551 : tab = 23'b11100110100010001100100;
12'd2552 : tab = 23'b11100110011100000110000;
12'd2553 : tab = 23'b11100110010101111111110;
12'd2554 : tab = 23'b11100110001111111001110;
12'd2555 : tab = 23'b11100110001001110100001;
12'd2556 : tab = 23'b11100110000011101110100;
12'd2557 : tab = 23'b11100101111101101001010;
12'd2558 : tab = 23'b11100101110111100100011;
12'd2559 : tab = 23'b11100101110001011111100;
12'd2560 : tab = 23'b11100101101011011011000;
12'd2561 : tab = 23'b11100101100101010110100;
12'd2562 : tab = 23'b11100101011111010010011;
12'd2563 : tab = 23'b11100101011001001110101;
12'd2564 : tab = 23'b11100101010011001010111;
12'd2565 : tab = 23'b11100101001101000111100;
12'd2566 : tab = 23'b11100101000111000100001;
12'd2567 : tab = 23'b11100101000001000001001;
12'd2568 : tab = 23'b11100100111010111110010;
12'd2569 : tab = 23'b11100100110100111011111;
12'd2570 : tab = 23'b11100100101110111001101;
12'd2571 : tab = 23'b11100100101000110111100;
12'd2572 : tab = 23'b11100100100010110101100;
12'd2573 : tab = 23'b11100100011100110100000;
12'd2574 : tab = 23'b11100100010110110010100;
12'd2575 : tab = 23'b11100100010000110001011;
12'd2576 : tab = 23'b11100100001010110000100;
12'd2577 : tab = 23'b11100100000100101111110;
12'd2578 : tab = 23'b11100011111110101111001;
12'd2579 : tab = 23'b11100011111000101110110;
12'd2580 : tab = 23'b11100011110010101110110;
12'd2581 : tab = 23'b11100011101100101111000;
12'd2582 : tab = 23'b11100011100110101111010;
12'd2583 : tab = 23'b11100011100000101111111;
12'd2584 : tab = 23'b11100011011010110000101;
12'd2585 : tab = 23'b11100011010100110001110;
12'd2586 : tab = 23'b11100011001110110011000;
12'd2587 : tab = 23'b11100011001000110100011;
12'd2588 : tab = 23'b11100011000010110110010;
12'd2589 : tab = 23'b11100010111100111000001;
12'd2590 : tab = 23'b11100010110110111010011;
12'd2591 : tab = 23'b11100010110000111100101;
12'd2592 : tab = 23'b11100010101010111111010;
12'd2593 : tab = 23'b11100010100101000010000;
12'd2594 : tab = 23'b11100010011111000101000;
12'd2595 : tab = 23'b11100010011001001000010;
12'd2596 : tab = 23'b11100010010011001011110;
12'd2597 : tab = 23'b11100010001101001111011;
12'd2598 : tab = 23'b11100010000111010011100;
12'd2599 : tab = 23'b11100010000001010111101;
12'd2600 : tab = 23'b11100001111011011100000;
12'd2601 : tab = 23'b11100001110101100000101;
12'd2602 : tab = 23'b11100001101111100101010;
12'd2603 : tab = 23'b11100001101001101010011;
12'd2604 : tab = 23'b11100001100011101111101;
12'd2605 : tab = 23'b11100001011101110101000;
12'd2606 : tab = 23'b11100001010111111010100;
12'd2607 : tab = 23'b11100001010010000000100;
12'd2608 : tab = 23'b11100001001100000110100;
12'd2609 : tab = 23'b11100001000110001100111;
12'd2610 : tab = 23'b11100001000000010011100;
12'd2611 : tab = 23'b11100000111010011010010;
12'd2612 : tab = 23'b11100000110100100001001;
12'd2613 : tab = 23'b11100000101110101000010;
12'd2614 : tab = 23'b11100000101000101111110;
12'd2615 : tab = 23'b11100000100010110111010;
12'd2616 : tab = 23'b11100000011100111111001;
12'd2617 : tab = 23'b11100000010111000111010;
12'd2618 : tab = 23'b11100000010001001111100;
12'd2619 : tab = 23'b11100000001011010111111;
12'd2620 : tab = 23'b11100000000101100000100;
12'd2621 : tab = 23'b11011111111111101001100;
12'd2622 : tab = 23'b11011111111001110010110;
12'd2623 : tab = 23'b11011111110011111011111;
12'd2624 : tab = 23'b11011111101110000101101;
12'd2625 : tab = 23'b11011111101000001111011;
12'd2626 : tab = 23'b11011111100010011001010;
12'd2627 : tab = 23'b11011111011100100011101;
12'd2628 : tab = 23'b11011111010110101110000;
12'd2629 : tab = 23'b11011111010000111000101;
12'd2630 : tab = 23'b11011111001011000011001;
12'd2631 : tab = 23'b11011111000101001110011;
12'd2632 : tab = 23'b11011110111111011001101;
12'd2633 : tab = 23'b11011110111001100101010;
12'd2634 : tab = 23'b11011110110011110000111;
12'd2635 : tab = 23'b11011110101101111100100;
12'd2636 : tab = 23'b11011110101000001000111;
12'd2637 : tab = 23'b11011110100010010101010;
12'd2638 : tab = 23'b11011110011100100001101;
12'd2639 : tab = 23'b11011110010110101110011;
12'd2640 : tab = 23'b11011110010000111011010;
12'd2641 : tab = 23'b11011110001011001000101;
12'd2642 : tab = 23'b11011110000101010101110;
12'd2643 : tab = 23'b11011101111111100011100;
12'd2644 : tab = 23'b11011101111001110001001;
12'd2645 : tab = 23'b11011101110011111111011;
12'd2646 : tab = 23'b11011101101110001101010;
12'd2647 : tab = 23'b11011101101000011011111;
12'd2648 : tab = 23'b11011101100010101010100;
12'd2649 : tab = 23'b11011101011100111001010;
12'd2650 : tab = 23'b11011101010111001000100;
12'd2651 : tab = 23'b11011101010001010111110;
12'd2652 : tab = 23'b11011101001011100111000;
12'd2653 : tab = 23'b11011101000101110110101;
12'd2654 : tab = 23'b11011101000000000110110;
12'd2655 : tab = 23'b11011100111010010110111;
12'd2656 : tab = 23'b11011100110100100111000;
12'd2657 : tab = 23'b11011100101110110111100;
12'd2658 : tab = 23'b11011100101001001000010;
12'd2659 : tab = 23'b11011100100011011001010;
12'd2660 : tab = 23'b11011100011101101010010;
12'd2661 : tab = 23'b11011100010111111011110;
12'd2662 : tab = 23'b11011100010010001101000;
12'd2663 : tab = 23'b11011100001100011110110;
12'd2664 : tab = 23'b11011100000110110000110;
12'd2665 : tab = 23'b11011100000001000011000;
12'd2666 : tab = 23'b11011011111011010101011;
12'd2667 : tab = 23'b11011011110101101000000;
12'd2668 : tab = 23'b11011011101111111010110;
12'd2669 : tab = 23'b11011011101010001101101;
12'd2670 : tab = 23'b11011011100100100000110;
12'd2671 : tab = 23'b11011011011110110100010;
12'd2672 : tab = 23'b11011011011001000111110;
12'd2673 : tab = 23'b11011011010011011011101;
12'd2674 : tab = 23'b11011011001101101111110;
12'd2675 : tab = 23'b11011011001000000011110;
12'd2676 : tab = 23'b11011011000010011000010;
12'd2677 : tab = 23'b11011010111100101100110;
12'd2678 : tab = 23'b11011010110111000001101;
12'd2679 : tab = 23'b11011010110001010110101;
12'd2680 : tab = 23'b11011010101011101100000;
12'd2681 : tab = 23'b11011010100110000001011;
12'd2682 : tab = 23'b11011010100000010111001;
12'd2683 : tab = 23'b11011010011010101100111;
12'd2684 : tab = 23'b11011010010101000011000;
12'd2685 : tab = 23'b11011010001111011001001;
12'd2686 : tab = 23'b11011010001001101111101;
12'd2687 : tab = 23'b11011010000100000110001;
12'd2688 : tab = 23'b11011001111110011101000;
12'd2689 : tab = 23'b11011001111000110100000;
12'd2690 : tab = 23'b11011001110011001011001;
12'd2691 : tab = 23'b11011001101101100010110;
12'd2692 : tab = 23'b11011001100111111010011;
12'd2693 : tab = 23'b11011001100010010010010;
12'd2694 : tab = 23'b11011001011100101010011;
12'd2695 : tab = 23'b11011001010111000010011;
12'd2696 : tab = 23'b11011001010001011011001;
12'd2697 : tab = 23'b11011001001011110011110;
12'd2698 : tab = 23'b11011001000110001100100;
12'd2699 : tab = 23'b11011001000000100101011;
12'd2700 : tab = 23'b11011000111010111110111;
12'd2701 : tab = 23'b11011000110101011000011;
12'd2702 : tab = 23'b11011000101111110001111;
12'd2703 : tab = 23'b11011000101010001011110;
12'd2704 : tab = 23'b11011000100100100101101;
12'd2705 : tab = 23'b11011000011110111111111;
12'd2706 : tab = 23'b11011000011001011010100;
12'd2707 : tab = 23'b11011000010011110101001;
12'd2708 : tab = 23'b11011000001110001111110;
12'd2709 : tab = 23'b11011000001000101011000;
12'd2710 : tab = 23'b11011000000011000110001;
12'd2711 : tab = 23'b11010111111101100001100;
12'd2712 : tab = 23'b11010111110111111101010;
12'd2713 : tab = 23'b11010111110010011001000;
12'd2714 : tab = 23'b11010111101100110101001;
12'd2715 : tab = 23'b11010111100111010001010;
12'd2716 : tab = 23'b11010111100001101101110;
12'd2717 : tab = 23'b11010111011100001010010;
12'd2718 : tab = 23'b11010111010110100111001;
12'd2719 : tab = 23'b11010111010001000100000;
12'd2720 : tab = 23'b11010111001011100001010;
12'd2721 : tab = 23'b11010111000101111110110;
12'd2722 : tab = 23'b11010111000000011100001;
12'd2723 : tab = 23'b11010110111010111010001;
12'd2724 : tab = 23'b11010110110101011000001;
12'd2725 : tab = 23'b11010110101111110110001;
12'd2726 : tab = 23'b11010110101010010100100;
12'd2727 : tab = 23'b11010110100100110011010;
12'd2728 : tab = 23'b11010110011111010010000;
12'd2729 : tab = 23'b11010110011001110000110;
12'd2730 : tab = 23'b11010110010100001111111;
12'd2731 : tab = 23'b11010110001110101111011;
12'd2732 : tab = 23'b11010110001001001110111;
12'd2733 : tab = 23'b11010110000011101110100;
12'd2734 : tab = 23'b11010101111110001110101;
12'd2735 : tab = 23'b11010101111000101110110;
12'd2736 : tab = 23'b11010101110011001111001;
12'd2737 : tab = 23'b11010101101101101111011;
12'd2738 : tab = 23'b11010101101000010000000;
12'd2739 : tab = 23'b11010101100010110001000;
12'd2740 : tab = 23'b11010101011101010010000;
12'd2741 : tab = 23'b11010101010111110011011;
12'd2742 : tab = 23'b11010101010010010100110;
12'd2743 : tab = 23'b11010101001100110110100;
12'd2744 : tab = 23'b11010101000111011000010;
12'd2745 : tab = 23'b11010101000001111010011;
12'd2746 : tab = 23'b11010100111100011100100;
12'd2747 : tab = 23'b11010100110110111111000;
12'd2748 : tab = 23'b11010100110001100001100;
12'd2749 : tab = 23'b11010100101100000100011;
12'd2750 : tab = 23'b11010100100110100111010;
12'd2751 : tab = 23'b11010100100001001010100;
12'd2752 : tab = 23'b11010100011011101101110;
12'd2753 : tab = 23'b11010100010110010001011;
12'd2754 : tab = 23'b11010100010000110101010;
12'd2755 : tab = 23'b11010100001011011001000;
12'd2756 : tab = 23'b11010100000101111101010;
12'd2757 : tab = 23'b11010100000000100001100;
12'd2758 : tab = 23'b11010011111011000110001;
12'd2759 : tab = 23'b11010011110101101010111;
12'd2760 : tab = 23'b11010011110000001111101;
12'd2761 : tab = 23'b11010011101010110100110;
12'd2762 : tab = 23'b11010011100101011001111;
12'd2763 : tab = 23'b11010011011111111111011;
12'd2764 : tab = 23'b11010011011010100101000;
12'd2765 : tab = 23'b11010011010101001010110;
12'd2766 : tab = 23'b11010011001111110001000;
12'd2767 : tab = 23'b11010011001010010111010;
12'd2768 : tab = 23'b11010011000100111101100;
12'd2769 : tab = 23'b11010010111111100100001;
12'd2770 : tab = 23'b11010010111010001010110;
12'd2771 : tab = 23'b11010010110100110001110;
12'd2772 : tab = 23'b11010010101111011000110;
12'd2773 : tab = 23'b11010010101010000000001;
12'd2774 : tab = 23'b11010010100100100111110;
12'd2775 : tab = 23'b11010010011111001111010;
12'd2776 : tab = 23'b11010010011001110111011;
12'd2777 : tab = 23'b11010010010100011111001;
12'd2778 : tab = 23'b11010010001111000111101;
12'd2779 : tab = 23'b11010010001001110000000;
12'd2780 : tab = 23'b11010010000100011000101;
12'd2781 : tab = 23'b11010001111111000001100;
12'd2782 : tab = 23'b11010001111001101010011;
12'd2783 : tab = 23'b11010001110100010011101;
12'd2784 : tab = 23'b11010001101110111100111;
12'd2785 : tab = 23'b11010001101001100110100;
12'd2786 : tab = 23'b11010001100100010000001;
12'd2787 : tab = 23'b11010001011110111010001;
12'd2788 : tab = 23'b11010001011001100100001;
12'd2789 : tab = 23'b11010001010100001110100;
12'd2790 : tab = 23'b11010001001110111000111;
12'd2791 : tab = 23'b11010001001001100011101;
12'd2792 : tab = 23'b11010001000100001110011;
12'd2793 : tab = 23'b11010000111110111001100;
12'd2794 : tab = 23'b11010000111001100100101;
12'd2795 : tab = 23'b11010000110100010000001;
12'd2796 : tab = 23'b11010000101110111011101;
12'd2797 : tab = 23'b11010000101001100111100;
12'd2798 : tab = 23'b11010000100100010011011;
12'd2799 : tab = 23'b11010000011110111111100;
12'd2800 : tab = 23'b11010000011001101011110;
12'd2801 : tab = 23'b11010000010100011000010;
12'd2802 : tab = 23'b11010000001111000100110;
12'd2803 : tab = 23'b11010000001001110001100;
12'd2804 : tab = 23'b11010000000100011110110;
12'd2805 : tab = 23'b11001111111111001100000;
12'd2806 : tab = 23'b11001111111001111001010;
12'd2807 : tab = 23'b11001111110100100110111;
12'd2808 : tab = 23'b11001111101111010100101;
12'd2809 : tab = 23'b11001111101010000010100;
12'd2810 : tab = 23'b11001111100100110000100;
12'd2811 : tab = 23'b11001111011111011111000;
12'd2812 : tab = 23'b11001111011010001101100;
12'd2813 : tab = 23'b11001111010100111100000;
12'd2814 : tab = 23'b11001111001111101010111;
12'd2815 : tab = 23'b11001111001010011001110;
12'd2816 : tab = 23'b11001111000101001001000;
12'd2817 : tab = 23'b11001110111111111000100;
12'd2818 : tab = 23'b11001110111010100111111;
12'd2819 : tab = 23'b11001110110101010111110;
12'd2820 : tab = 23'b11001110110000000111100;
12'd2821 : tab = 23'b11001110101010110111100;
12'd2822 : tab = 23'b11001110100101100111111;
12'd2823 : tab = 23'b11001110100000011000010;
12'd2824 : tab = 23'b11001110011011001001000;
12'd2825 : tab = 23'b11001110010101111001110;
12'd2826 : tab = 23'b11001110010000101010110;
12'd2827 : tab = 23'b11001110001011011100000;
12'd2828 : tab = 23'b11001110000110001101001;
12'd2829 : tab = 23'b11001110000000111110101;
12'd2830 : tab = 23'b11001101111011110000100;
12'd2831 : tab = 23'b11001101110110100010010;
12'd2832 : tab = 23'b11001101110001010100010;
12'd2833 : tab = 23'b11001101101100000110100;
12'd2834 : tab = 23'b11001101100110111000110;
12'd2835 : tab = 23'b11001101100001101011011;
12'd2836 : tab = 23'b11001101011100011110010;
12'd2837 : tab = 23'b11001101010111010001000;
12'd2838 : tab = 23'b11001101010010000100011;
12'd2839 : tab = 23'b11001101001100110111011;
12'd2840 : tab = 23'b11001101000111101010110;
12'd2841 : tab = 23'b11001101000010011110100;
12'd2842 : tab = 23'b11001100111101010010010;
12'd2843 : tab = 23'b11001100111000000110011;
12'd2844 : tab = 23'b11001100110010111010100;
12'd2845 : tab = 23'b11001100101101101110101;
12'd2846 : tab = 23'b11001100101000100011001;
12'd2847 : tab = 23'b11001100100011011000000;
12'd2848 : tab = 23'b11001100011110001100111;
12'd2849 : tab = 23'b11001100011001000001110;
12'd2850 : tab = 23'b11001100010011110111000;
12'd2851 : tab = 23'b11001100001110101100010;
12'd2852 : tab = 23'b11001100001001100001111;
12'd2853 : tab = 23'b11001100000100010111100;
12'd2854 : tab = 23'b11001011111111001101100;
12'd2855 : tab = 23'b11001011111010000011100;
12'd2856 : tab = 23'b11001011110100111001111;
12'd2857 : tab = 23'b11001011101111110000010;
12'd2858 : tab = 23'b11001011101010100110110;
12'd2859 : tab = 23'b11001011100101011101100;
12'd2860 : tab = 23'b11001011100000010100100;
12'd2861 : tab = 23'b11001011011011001011101;
12'd2862 : tab = 23'b11001011010110000010110;
12'd2863 : tab = 23'b11001011010000111010010;
12'd2864 : tab = 23'b11001011001011110010000;
12'd2865 : tab = 23'b11001011000110101001101;
12'd2866 : tab = 23'b11001011000001100001100;
12'd2867 : tab = 23'b11001010111100011001110;
12'd2868 : tab = 23'b11001010110111010010000;
12'd2869 : tab = 23'b11001010110010001010101;
12'd2870 : tab = 23'b11001010101101000011010;
12'd2871 : tab = 23'b11001010100111111100000;
12'd2872 : tab = 23'b11001010100010110100111;
12'd2873 : tab = 23'b11001010011101101110010;
12'd2874 : tab = 23'b11001010011000100111101;
12'd2875 : tab = 23'b11001010010011100001000;
12'd2876 : tab = 23'b11001010001110011010110;
12'd2877 : tab = 23'b11001010001001010100100;
12'd2878 : tab = 23'b11001010000100001110101;
12'd2879 : tab = 23'b11001001111111001000110;
12'd2880 : tab = 23'b11001001111010000011000;
12'd2881 : tab = 23'b11001001110100111101100;
12'd2882 : tab = 23'b11001001101111111000010;
12'd2883 : tab = 23'b11001001101010110011001;
12'd2884 : tab = 23'b11001001100101101110010;
12'd2885 : tab = 23'b11001001100000101001010;
12'd2886 : tab = 23'b11001001011011100100110;
12'd2887 : tab = 23'b11001001010110100000001;
12'd2888 : tab = 23'b11001001010001011011110;
12'd2889 : tab = 23'b11001001001100010111110;
12'd2890 : tab = 23'b11001001000111010011110;
12'd2891 : tab = 23'b11001001000010010000000;
12'd2892 : tab = 23'b11001000111101001100100;
12'd2893 : tab = 23'b11001000111000001000111;
12'd2894 : tab = 23'b11001000110011000101101;
12'd2895 : tab = 23'b11001000101110000010011;
12'd2896 : tab = 23'b11001000101000111111100;
12'd2897 : tab = 23'b11001000100011111100110;
12'd2898 : tab = 23'b11001000011110111010001;
12'd2899 : tab = 23'b11001000011001110111101;
12'd2900 : tab = 23'b11001000010100110101100;
12'd2901 : tab = 23'b11001000001111110011011;
12'd2902 : tab = 23'b11001000001010110001010;
12'd2903 : tab = 23'b11001000000101101111100;
12'd2904 : tab = 23'b11001000000000101110000;
12'd2905 : tab = 23'b11000111111011101100011;
12'd2906 : tab = 23'b11000111110110101011010;
12'd2907 : tab = 23'b11000111110001101010000;
12'd2908 : tab = 23'b11000111101100101001000;
12'd2909 : tab = 23'b11000111100111101000011;
12'd2910 : tab = 23'b11000111100010100111110;
12'd2911 : tab = 23'b11000111011101100111001;
12'd2912 : tab = 23'b11000111011000100110111;
12'd2913 : tab = 23'b11000111010011100110110;
12'd2914 : tab = 23'b11000111001110100110110;
12'd2915 : tab = 23'b11000111001001100111000;
12'd2916 : tab = 23'b11000111000100100111011;
12'd2917 : tab = 23'b11000110111111100111111;
12'd2918 : tab = 23'b11000110111010101000100;
12'd2919 : tab = 23'b11000110110101101001100;
12'd2920 : tab = 23'b11000110110000101010100;
12'd2921 : tab = 23'b11000110101011101011110;
12'd2922 : tab = 23'b11000110100110101101000;
12'd2923 : tab = 23'b11000110100001101110101;
12'd2924 : tab = 23'b11000110011100110000010;
12'd2925 : tab = 23'b11000110010111110001111;
12'd2926 : tab = 23'b11000110010010110011111;
12'd2927 : tab = 23'b11000110001101110110000;
12'd2928 : tab = 23'b11000110001000111000100;
12'd2929 : tab = 23'b11000110000011111011000;
12'd2930 : tab = 23'b11000101111110111101100;
12'd2931 : tab = 23'b11000101111010000000100;
12'd2932 : tab = 23'b11000101110101000011100;
12'd2933 : tab = 23'b11000101110000000110100;
12'd2934 : tab = 23'b11000101101011001001111;
12'd2935 : tab = 23'b11000101100110001101011;
12'd2936 : tab = 23'b11000101100001010000111;
12'd2937 : tab = 23'b11000101011100010100110;
12'd2938 : tab = 23'b11000101010111011000101;
12'd2939 : tab = 23'b11000101010010011100111;
12'd2940 : tab = 23'b11000101001101100001001;
12'd2941 : tab = 23'b11000101001000100101011;
12'd2942 : tab = 23'b11000101000011101010000;
12'd2943 : tab = 23'b11000100111110101110110;
12'd2944 : tab = 23'b11000100111001110011101;
12'd2945 : tab = 23'b11000100110100111000101;
12'd2946 : tab = 23'b11000100101111111110000;
12'd2947 : tab = 23'b11000100101011000011011;
12'd2948 : tab = 23'b11000100100110001001000;
12'd2949 : tab = 23'b11000100100001001110110;
12'd2950 : tab = 23'b11000100011100010100100;
12'd2951 : tab = 23'b11000100010111011010100;
12'd2952 : tab = 23'b11000100010010100000111;
12'd2953 : tab = 23'b11000100001101100111000;
12'd2954 : tab = 23'b11000100001000101101100;
12'd2955 : tab = 23'b11000100000011110100010;
12'd2956 : tab = 23'b11000011111110111011000;
12'd2957 : tab = 23'b11000011111010000010001;
12'd2958 : tab = 23'b11000011110101001001010;
12'd2959 : tab = 23'b11000011110000010000101;
12'd2960 : tab = 23'b11000011101011010111111;
12'd2961 : tab = 23'b11000011100110011111110;
12'd2962 : tab = 23'b11000011100001100111100;
12'd2963 : tab = 23'b11000011011100101111010;
12'd2964 : tab = 23'b11000011010111110111100;
12'd2965 : tab = 23'b11000011010010111111110;
12'd2966 : tab = 23'b11000011001110001000010;
12'd2967 : tab = 23'b11000011001001010000101;
12'd2968 : tab = 23'b11000011000100011001011;
12'd2969 : tab = 23'b11000010111111100010010;
12'd2970 : tab = 23'b11000010111010101011010;
12'd2971 : tab = 23'b11000010110101110100011;
12'd2972 : tab = 23'b11000010110000111101111;
12'd2973 : tab = 23'b11000010101100000111011;
12'd2974 : tab = 23'b11000010100111010000111;
12'd2975 : tab = 23'b11000010100010011010110;
12'd2976 : tab = 23'b11000010011101100100110;
12'd2977 : tab = 23'b11000010011000101110111;
12'd2978 : tab = 23'b11000010010011111001001;
12'd2979 : tab = 23'b11000010001111000011110;
12'd2980 : tab = 23'b11000010001010001110011;
12'd2981 : tab = 23'b11000010000101011001000;
12'd2982 : tab = 23'b11000010000000100100000;
12'd2983 : tab = 23'b11000001111011101111000;
12'd2984 : tab = 23'b11000001110110111010011;
12'd2985 : tab = 23'b11000001110010000101110;
12'd2986 : tab = 23'b11000001101101010001001;
12'd2987 : tab = 23'b11000001101000011100111;
12'd2988 : tab = 23'b11000001100011101000101;
12'd2989 : tab = 23'b11000001011110110100110;
12'd2990 : tab = 23'b11000001011010000000111;
12'd2991 : tab = 23'b11000001010101001101000;
12'd2992 : tab = 23'b11000001010000011001100;
12'd2993 : tab = 23'b11000001001011100110011;
12'd2994 : tab = 23'b11000001000110110010111;
12'd2995 : tab = 23'b11000001000010000000000;
12'd2996 : tab = 23'b11000000111101001101000;
12'd2997 : tab = 23'b11000000111000011010010;
12'd2998 : tab = 23'b11000000110011100111110;
12'd2999 : tab = 23'b11000000101110110101001;
12'd3000 : tab = 23'b11000000101010000010110;
12'd3001 : tab = 23'b11000000100101010000110;
12'd3002 : tab = 23'b11000000100000011110110;
12'd3003 : tab = 23'b11000000011011101100110;
12'd3004 : tab = 23'b11000000010110111011001;
12'd3005 : tab = 23'b11000000010010001001100;
12'd3006 : tab = 23'b11000000001101011000010;
12'd3007 : tab = 23'b11000000001000100111000;
12'd3008 : tab = 23'b11000000000011110101110;
12'd3009 : tab = 23'b10111111111111000100111;
12'd3010 : tab = 23'b10111111111010010100000;
12'd3011 : tab = 23'b10111111110101100011100;
12'd3012 : tab = 23'b10111111110000110011000;
12'd3013 : tab = 23'b10111111101100000010110;
12'd3014 : tab = 23'b10111111100111010010011;
12'd3015 : tab = 23'b10111111100010100010101;
12'd3016 : tab = 23'b10111111011101110010110;
12'd3017 : tab = 23'b10111111011001000011000;
12'd3018 : tab = 23'b10111111010100010011011;
12'd3019 : tab = 23'b10111111001111100100000;
12'd3020 : tab = 23'b10111111001010110100101;
12'd3021 : tab = 23'b10111111000110000101101;
12'd3022 : tab = 23'b10111111000001010110101;
12'd3023 : tab = 23'b10111110111100100111110;
12'd3024 : tab = 23'b10111110110111111001000;
12'd3025 : tab = 23'b10111110110011001010100;
12'd3026 : tab = 23'b10111110101110011100001;
12'd3027 : tab = 23'b10111110101001101101111;
12'd3028 : tab = 23'b10111110100100111111110;
12'd3029 : tab = 23'b10111110100000010010001;
12'd3030 : tab = 23'b10111110011011100100010;
12'd3031 : tab = 23'b10111110010110110110100;
12'd3032 : tab = 23'b10111110010010001001010;
12'd3033 : tab = 23'b10111110001101011011110;
12'd3034 : tab = 23'b10111110001000101110101;
12'd3035 : tab = 23'b10111110000100000001100;
12'd3036 : tab = 23'b10111101111111010100110;
12'd3037 : tab = 23'b10111101111010101000000;
12'd3038 : tab = 23'b10111101110101111011010;
12'd3039 : tab = 23'b10111101110001001110111;
12'd3040 : tab = 23'b10111101101100100010110;
12'd3041 : tab = 23'b10111101100111110110100;
12'd3042 : tab = 23'b10111101100011001010100;
12'd3043 : tab = 23'b10111101011110011110110;
12'd3044 : tab = 23'b10111101011001110010111;
12'd3045 : tab = 23'b10111101010101000111101;
12'd3046 : tab = 23'b10111101010000011100010;
12'd3047 : tab = 23'b10111101001011110000110;
12'd3048 : tab = 23'b10111101000111000101111;
12'd3049 : tab = 23'b10111101000010011010110;
12'd3050 : tab = 23'b10111100111101110000000;
12'd3051 : tab = 23'b10111100111001000101010;
12'd3052 : tab = 23'b10111100110100011010110;
12'd3053 : tab = 23'b10111100101111110000100;
12'd3054 : tab = 23'b10111100101011000110001;
12'd3055 : tab = 23'b10111100100110011100010;
12'd3056 : tab = 23'b10111100100001110010010;
12'd3057 : tab = 23'b10111100011101001000100;
12'd3058 : tab = 23'b10111100011000011110110;
12'd3059 : tab = 23'b10111100010011110101011;
12'd3060 : tab = 23'b10111100001111001100000;
12'd3061 : tab = 23'b10111100001010100010110;
12'd3062 : tab = 23'b10111100000101111001101;
12'd3063 : tab = 23'b10111100000001010000110;
12'd3064 : tab = 23'b10111011111100101000000;
12'd3065 : tab = 23'b10111011110111111111011;
12'd3066 : tab = 23'b10111011110011010111001;
12'd3067 : tab = 23'b10111011101110101110110;
12'd3068 : tab = 23'b10111011101010000110100;
12'd3069 : tab = 23'b10111011100101011110011;
12'd3070 : tab = 23'b10111011100000110110100;
12'd3071 : tab = 23'b10111011011100001110101;
12'd3072 : tab = 23'b10111011010111100111001;
12'd3073 : tab = 23'b10111011010010111111101;
12'd3074 : tab = 23'b10111011001110011000100;
12'd3075 : tab = 23'b10111011001001110001010;
12'd3076 : tab = 23'b10111011000101001010010;
12'd3077 : tab = 23'b10111011000000100011010;
12'd3078 : tab = 23'b10111010111011111100110;
12'd3079 : tab = 23'b10111010110111010110000;
12'd3080 : tab = 23'b10111010110010101111100;
12'd3081 : tab = 23'b10111010101110001001010;
12'd3082 : tab = 23'b10111010101001100011000;
12'd3083 : tab = 23'b10111010100100111101000;
12'd3084 : tab = 23'b10111010100000010111000;
12'd3085 : tab = 23'b10111010011011110001100;
12'd3086 : tab = 23'b10111010010111001011110;
12'd3087 : tab = 23'b10111010010010100110011;
12'd3088 : tab = 23'b10111010001110000001001;
12'd3089 : tab = 23'b10111010001001011011111;
12'd3090 : tab = 23'b10111010000100110110110;
12'd3091 : tab = 23'b10111010000000010010001;
12'd3092 : tab = 23'b10111001111011101101010;
12'd3093 : tab = 23'b10111001110111001000110;
12'd3094 : tab = 23'b10111001110010100100010;
12'd3095 : tab = 23'b10111001101110000000000;
12'd3096 : tab = 23'b10111001101001011011101;
12'd3097 : tab = 23'b10111001100100110111100;
12'd3098 : tab = 23'b10111001100000010011110;
12'd3099 : tab = 23'b10111001011011110000000;
12'd3100 : tab = 23'b10111001010111001100010;
12'd3101 : tab = 23'b10111001010010101000111;
12'd3102 : tab = 23'b10111001001110000101100;
12'd3103 : tab = 23'b10111001001001100010100;
12'd3104 : tab = 23'b10111001000100111111010;
12'd3105 : tab = 23'b10111001000000011100100;
12'd3106 : tab = 23'b10111000111011111001110;
12'd3107 : tab = 23'b10111000110111010111010;
12'd3108 : tab = 23'b10111000110010110100101;
12'd3109 : tab = 23'b10111000101110010010011;
12'd3110 : tab = 23'b10111000101001110000001;
12'd3111 : tab = 23'b10111000100101001110000;
12'd3112 : tab = 23'b10111000100000101100010;
12'd3113 : tab = 23'b10111000011100001010010;
12'd3114 : tab = 23'b10111000010111101000101;
12'd3115 : tab = 23'b10111000010011000111001;
12'd3116 : tab = 23'b10111000001110100101110;
12'd3117 : tab = 23'b10111000001010000100100;
12'd3118 : tab = 23'b10111000000101100011011;
12'd3119 : tab = 23'b10111000000001000010101;
12'd3120 : tab = 23'b10110111111100100001110;
12'd3121 : tab = 23'b10110111111000000001001;
12'd3122 : tab = 23'b10110111110011100000100;
12'd3123 : tab = 23'b10110111101111000000010;
12'd3124 : tab = 23'b10110111101010100000000;
12'd3125 : tab = 23'b10110111100101111111110;
12'd3126 : tab = 23'b10110111100001011111110;
12'd3127 : tab = 23'b10110111011101000000000;
12'd3128 : tab = 23'b10110111011000100000011;
12'd3129 : tab = 23'b10110111010100000000110;
12'd3130 : tab = 23'b10110111001111100001010;
12'd3131 : tab = 23'b10110111001011000010000;
12'd3132 : tab = 23'b10110111000110100010110;
12'd3133 : tab = 23'b10110111000010000011110;
12'd3134 : tab = 23'b10110110111101100100111;
12'd3135 : tab = 23'b10110110111001000110011;
12'd3136 : tab = 23'b10110110110100100111110;
12'd3137 : tab = 23'b10110110110000001001010;
12'd3138 : tab = 23'b10110110101011101010111;
12'd3139 : tab = 23'b10110110100111001100100;
12'd3140 : tab = 23'b10110110100010101110101;
12'd3141 : tab = 23'b10110110011110010000110;
12'd3142 : tab = 23'b10110110011001110010110;
12'd3143 : tab = 23'b10110110010101010101011;
12'd3144 : tab = 23'b10110110010000110111101;
12'd3145 : tab = 23'b10110110001100011010010;
12'd3146 : tab = 23'b10110110000111111101010;
12'd3147 : tab = 23'b10110110000011100000000;
12'd3148 : tab = 23'b10110101111111000011010;
12'd3149 : tab = 23'b10110101111010100110010;
12'd3150 : tab = 23'b10110101110110001001101;
12'd3151 : tab = 23'b10110101110001101101000;
12'd3152 : tab = 23'b10110101101101010000100;
12'd3153 : tab = 23'b10110101101000110100010;
12'd3154 : tab = 23'b10110101100100011000010;
12'd3155 : tab = 23'b10110101011111111100000;
12'd3156 : tab = 23'b10110101011011100000001;
12'd3157 : tab = 23'b10110101010111000100101;
12'd3158 : tab = 23'b10110101010010101000110;
12'd3159 : tab = 23'b10110101001110001101010;
12'd3160 : tab = 23'b10110101001001110010001;
12'd3161 : tab = 23'b10110101000101010110110;
12'd3162 : tab = 23'b10110101000000111011111;
12'd3163 : tab = 23'b10110100111100100000110;
12'd3164 : tab = 23'b10110100111000000110000;
12'd3165 : tab = 23'b10110100110011101011100;
12'd3166 : tab = 23'b10110100101111010000111;
12'd3167 : tab = 23'b10110100101010110110100;
12'd3168 : tab = 23'b10110100100110011100001;
12'd3169 : tab = 23'b10110100100010000010001;
12'd3170 : tab = 23'b10110100011101101000001;
12'd3171 : tab = 23'b10110100011001001110001;
12'd3172 : tab = 23'b10110100010100110100100;
12'd3173 : tab = 23'b10110100010000011010111;
12'd3174 : tab = 23'b10110100001100000001010;
12'd3175 : tab = 23'b10110100000111101000000;
12'd3176 : tab = 23'b10110100000011001110110;
12'd3177 : tab = 23'b10110011111110110101110;
12'd3178 : tab = 23'b10110011111010011100110;
12'd3179 : tab = 23'b10110011110110000100001;
12'd3180 : tab = 23'b10110011110001101011010;
12'd3181 : tab = 23'b10110011101101010010110;
12'd3182 : tab = 23'b10110011101000111010010;
12'd3183 : tab = 23'b10110011100100100010001;
12'd3184 : tab = 23'b10110011100000001010000;
12'd3185 : tab = 23'b10110011011011110001111;
12'd3186 : tab = 23'b10110011010111011010001;
12'd3187 : tab = 23'b10110011010011000010011;
12'd3188 : tab = 23'b10110011001110101010101;
12'd3189 : tab = 23'b10110011001010010011010;
12'd3190 : tab = 23'b10110011000101111011111;
12'd3191 : tab = 23'b10110011000001100100110;
12'd3192 : tab = 23'b10110010111101001101100;
12'd3193 : tab = 23'b10110010111000110110100;
12'd3194 : tab = 23'b10110010110100011111111;
12'd3195 : tab = 23'b10110010110000001001000;
12'd3196 : tab = 23'b10110010101011110010101;
12'd3197 : tab = 23'b10110010100111011100000;
12'd3198 : tab = 23'b10110010100011000101110;
12'd3199 : tab = 23'b10110010011110101111100;
12'd3200 : tab = 23'b10110010011010011001101;
12'd3201 : tab = 23'b10110010010110000011100;
12'd3202 : tab = 23'b10110010010001101101111;
12'd3203 : tab = 23'b10110010001101011000010;
12'd3204 : tab = 23'b10110010001001000010110;
12'd3205 : tab = 23'b10110010000100101101011;
12'd3206 : tab = 23'b10110010000000010111111;
12'd3207 : tab = 23'b10110001111100000010110;
12'd3208 : tab = 23'b10110001110111101101110;
12'd3209 : tab = 23'b10110001110011011000111;
12'd3210 : tab = 23'b10110001101111000100001;
12'd3211 : tab = 23'b10110001101010101111100;
12'd3212 : tab = 23'b10110001100110011011000;
12'd3213 : tab = 23'b10110001100010000110101;
12'd3214 : tab = 23'b10110001011101110010101;
12'd3215 : tab = 23'b10110001011001011110100;
12'd3216 : tab = 23'b10110001010101001010010;
12'd3217 : tab = 23'b10110001010000110110101;
12'd3218 : tab = 23'b10110001001100100011000;
12'd3219 : tab = 23'b10110001001000001111011;
12'd3220 : tab = 23'b10110001000011111011110;
12'd3221 : tab = 23'b10110000111111101000100;
12'd3222 : tab = 23'b10110000111011010101010;
12'd3223 : tab = 23'b10110000110111000010010;
12'd3224 : tab = 23'b10110000110010101111010;
12'd3225 : tab = 23'b10110000101110011100100;
12'd3226 : tab = 23'b10110000101010001001110;
12'd3227 : tab = 23'b10110000100101110111010;
12'd3228 : tab = 23'b10110000100001100100110;
12'd3229 : tab = 23'b10110000011101010010100;
12'd3230 : tab = 23'b10110000011001000000010;
12'd3231 : tab = 23'b10110000010100101110010;
12'd3232 : tab = 23'b10110000010000011100010;
12'd3233 : tab = 23'b10110000001100001010100;
12'd3234 : tab = 23'b10110000000111111000110;
12'd3235 : tab = 23'b10110000000011100111011;
12'd3236 : tab = 23'b10101111111111010101110;
12'd3237 : tab = 23'b10101111111011000100101;
12'd3238 : tab = 23'b10101111110110110011010;
12'd3239 : tab = 23'b10101111110010100010010;
12'd3240 : tab = 23'b10101111101110010001101;
12'd3241 : tab = 23'b10101111101010000000101;
12'd3242 : tab = 23'b10101111100101110000000;
12'd3243 : tab = 23'b10101111100001011111011;
12'd3244 : tab = 23'b10101111011101001111001;
12'd3245 : tab = 23'b10101111011000111110111;
12'd3246 : tab = 23'b10101111010100101110101;
12'd3247 : tab = 23'b10101111010000011110100;
12'd3248 : tab = 23'b10101111001100001110111;
12'd3249 : tab = 23'b10101111000111111111000;
12'd3250 : tab = 23'b10101111000011101111001;
12'd3251 : tab = 23'b10101110111111011111101;
12'd3252 : tab = 23'b10101110111011010000001;
12'd3253 : tab = 23'b10101110110111000001000;
12'd3254 : tab = 23'b10101110110010110001111;
12'd3255 : tab = 23'b10101110101110100010110;
12'd3256 : tab = 23'b10101110101010010100000;
12'd3257 : tab = 23'b10101110100110000101010;
12'd3258 : tab = 23'b10101110100001110110100;
12'd3259 : tab = 23'b10101110011101101000001;
12'd3260 : tab = 23'b10101110011001011001110;
12'd3261 : tab = 23'b10101110010101001011011;
12'd3262 : tab = 23'b10101110010000111101010;
12'd3263 : tab = 23'b10101110001100101111000;
12'd3264 : tab = 23'b10101110001000100001011;
12'd3265 : tab = 23'b10101110000100010011011;
12'd3266 : tab = 23'b10101110000000000101110;
12'd3267 : tab = 23'b10101101111011111000001;
12'd3268 : tab = 23'b10101101110111101010111;
12'd3269 : tab = 23'b10101101110011011101101;
12'd3270 : tab = 23'b10101101101111010000011;
12'd3271 : tab = 23'b10101101101011000011010;
12'd3272 : tab = 23'b10101101100110110110100;
12'd3273 : tab = 23'b10101101100010101001110;
12'd3274 : tab = 23'b10101101011110011100111;
12'd3275 : tab = 23'b10101101011010010000011;
12'd3276 : tab = 23'b10101101010110000011111;
12'd3277 : tab = 23'b10101101010001110111110;
12'd3278 : tab = 23'b10101101001101101011101;
12'd3279 : tab = 23'b10101101001001011111100;
12'd3280 : tab = 23'b10101101000101010011011;
12'd3281 : tab = 23'b10101101000001000111101;
12'd3282 : tab = 23'b10101100111100111011111;
12'd3283 : tab = 23'b10101100111000110000100;
12'd3284 : tab = 23'b10101100110100100101000;
12'd3285 : tab = 23'b10101100110000011001110;
12'd3286 : tab = 23'b10101100101100001110011;
12'd3287 : tab = 23'b10101100101000000011011;
12'd3288 : tab = 23'b10101100100011111000011;
12'd3289 : tab = 23'b10101100011111101101100;
12'd3290 : tab = 23'b10101100011011100010110;
12'd3291 : tab = 23'b10101100010111011000001;
12'd3292 : tab = 23'b10101100010011001101111;
12'd3293 : tab = 23'b10101100001111000011100;
12'd3294 : tab = 23'b10101100001010111001011;
12'd3295 : tab = 23'b10101100000110101111001;
12'd3296 : tab = 23'b10101100000010100101000;
12'd3297 : tab = 23'b10101011111110011011010;
12'd3298 : tab = 23'b10101011111010010001100;
12'd3299 : tab = 23'b10101011110110001000000;
12'd3300 : tab = 23'b10101011110001111110100;
12'd3301 : tab = 23'b10101011101101110101000;
12'd3302 : tab = 23'b10101011101001101011110;
12'd3303 : tab = 23'b10101011100101100010100;
12'd3304 : tab = 23'b10101011100001011001101;
12'd3305 : tab = 23'b10101011011101010000110;
12'd3306 : tab = 23'b10101011011001001000000;
12'd3307 : tab = 23'b10101011010100111111010;
12'd3308 : tab = 23'b10101011010000110110101;
12'd3309 : tab = 23'b10101011001100101110010;
12'd3310 : tab = 23'b10101011001000100101111;
12'd3311 : tab = 23'b10101011000100011101110;
12'd3312 : tab = 23'b10101011000000010101110;
12'd3313 : tab = 23'b10101010111100001101111;
12'd3314 : tab = 23'b10101010111000000101111;
12'd3315 : tab = 23'b10101010110011111110010;
12'd3316 : tab = 23'b10101010101111110110101;
12'd3317 : tab = 23'b10101010101011101111010;
12'd3318 : tab = 23'b10101010100111100111110;
12'd3319 : tab = 23'b10101010100011100000100;
12'd3320 : tab = 23'b10101010011111011001101;
12'd3321 : tab = 23'b10101010011011010010100;
12'd3322 : tab = 23'b10101010010111001011100;
12'd3323 : tab = 23'b10101010010011000101000;
12'd3324 : tab = 23'b10101010001110111110010;
12'd3325 : tab = 23'b10101010001010110111110;
12'd3326 : tab = 23'b10101010000110110001100;
12'd3327 : tab = 23'b10101010000010101011000;
12'd3328 : tab = 23'b10101001111110100100111;
12'd3329 : tab = 23'b10101001111010011110110;
12'd3330 : tab = 23'b10101001110110011001000;
12'd3331 : tab = 23'b10101001110010010011010;
12'd3332 : tab = 23'b10101001101110001101100;
12'd3333 : tab = 23'b10101001101010000111110;
12'd3334 : tab = 23'b10101001100110000010011;
12'd3335 : tab = 23'b10101001100001111101000;
12'd3336 : tab = 23'b10101001011101110111110;
12'd3337 : tab = 23'b10101001011001110010110;
12'd3338 : tab = 23'b10101001010101101101101;
12'd3339 : tab = 23'b10101001010001101001000;
12'd3340 : tab = 23'b10101001001101100100010;
12'd3341 : tab = 23'b10101001001001011111100;
12'd3342 : tab = 23'b10101001000101011011001;
12'd3343 : tab = 23'b10101001000001010110110;
12'd3344 : tab = 23'b10101000111101010010100;
12'd3345 : tab = 23'b10101000111001001110010;
12'd3346 : tab = 23'b10101000110101001010001;
12'd3347 : tab = 23'b10101000110001000110010;
12'd3348 : tab = 23'b10101000101101000010011;
12'd3349 : tab = 23'b10101000101000111110110;
12'd3350 : tab = 23'b10101000100100111011010;
12'd3351 : tab = 23'b10101000100000110111110;
12'd3352 : tab = 23'b10101000011100110100011;
12'd3353 : tab = 23'b10101000011000110001000;
12'd3354 : tab = 23'b10101000010100101110001;
12'd3355 : tab = 23'b10101000010000101011000;
12'd3356 : tab = 23'b10101000001100101000000;
12'd3357 : tab = 23'b10101000001000100101010;
12'd3358 : tab = 23'b10101000000100100010110;
12'd3359 : tab = 23'b10101000000000100000010;
12'd3360 : tab = 23'b10100111111100011101101;
12'd3361 : tab = 23'b10100111111000011011010;
12'd3362 : tab = 23'b10100111110100011001010;
12'd3363 : tab = 23'b10100111110000010111010;
12'd3364 : tab = 23'b10100111101100010101010;
12'd3365 : tab = 23'b10100111101000010011010;
12'd3366 : tab = 23'b10100111100100010001101;
12'd3367 : tab = 23'b10100111100000010000000;
12'd3368 : tab = 23'b10100111011100001110011;
12'd3369 : tab = 23'b10100111011000001101001;
12'd3370 : tab = 23'b10100111010100001011111;
12'd3371 : tab = 23'b10100111010000001010101;
12'd3372 : tab = 23'b10100111001100001001100;
12'd3373 : tab = 23'b10100111001000001000110;
12'd3374 : tab = 23'b10100111000100000111110;
12'd3375 : tab = 23'b10100111000000000111001;
12'd3376 : tab = 23'b10100110111100000110101;
12'd3377 : tab = 23'b10100110111000000110001;
12'd3378 : tab = 23'b10100110110100000101101;
12'd3379 : tab = 23'b10100110110000000101100;
12'd3380 : tab = 23'b10100110101100000101011;
12'd3381 : tab = 23'b10100110101000000101010;
12'd3382 : tab = 23'b10100110100100000101100;
12'd3383 : tab = 23'b10100110100000000101100;
12'd3384 : tab = 23'b10100110011100000110000;
12'd3385 : tab = 23'b10100110011000000110100;
12'd3386 : tab = 23'b10100110010100000110111;
12'd3387 : tab = 23'b10100110010000000111100;
12'd3388 : tab = 23'b10100110001100001000100;
12'd3389 : tab = 23'b10100110001000001001001;
12'd3390 : tab = 23'b10100110000100001010001;
12'd3391 : tab = 23'b10100110000000001011100;
12'd3392 : tab = 23'b10100101111100001100100;
12'd3393 : tab = 23'b10100101111000001101111;
12'd3394 : tab = 23'b10100101110100001111010;
12'd3395 : tab = 23'b10100101110000010001000;
12'd3396 : tab = 23'b10100101101100010010100;
12'd3397 : tab = 23'b10100101101000010100010;
12'd3398 : tab = 23'b10100101100100010110010;
12'd3399 : tab = 23'b10100101100000011000011;
12'd3400 : tab = 23'b10100101011100011010100;
12'd3401 : tab = 23'b10100101011000011100101;
12'd3402 : tab = 23'b10100101010100011111000;
12'd3403 : tab = 23'b10100101010000100001100;
12'd3404 : tab = 23'b10100101001100100100001;
12'd3405 : tab = 23'b10100101001000100110101;
12'd3406 : tab = 23'b10100101000100101001100;
12'd3407 : tab = 23'b10100101000000101100011;
12'd3408 : tab = 23'b10100100111100101111100;
12'd3409 : tab = 23'b10100100111000110010100;
12'd3410 : tab = 23'b10100100110100110101110;
12'd3411 : tab = 23'b10100100110000111001000;
12'd3412 : tab = 23'b10100100101100111100101;
12'd3413 : tab = 23'b10100100101001000000010;
12'd3414 : tab = 23'b10100100100101000011111;
12'd3415 : tab = 23'b10100100100001000111100;
12'd3416 : tab = 23'b10100100011101001011100;
12'd3417 : tab = 23'b10100100011001001111100;
12'd3418 : tab = 23'b10100100010101010011110;
12'd3419 : tab = 23'b10100100010001010111111;
12'd3420 : tab = 23'b10100100001101011100010;
12'd3421 : tab = 23'b10100100001001100000101;
12'd3422 : tab = 23'b10100100000101100101011;
12'd3423 : tab = 23'b10100100000001101010000;
12'd3424 : tab = 23'b10100011111101101110111;
12'd3425 : tab = 23'b10100011111001110011101;
12'd3426 : tab = 23'b10100011110101111000110;
12'd3427 : tab = 23'b10100011110001111101111;
12'd3428 : tab = 23'b10100011101110000011000;
12'd3429 : tab = 23'b10100011101010001000010;
12'd3430 : tab = 23'b10100011100110001101110;
12'd3431 : tab = 23'b10100011100010010011100;
12'd3432 : tab = 23'b10100011011110011001000;
12'd3433 : tab = 23'b10100011011010011110111;
12'd3434 : tab = 23'b10100011010110100100110;
12'd3435 : tab = 23'b10100011010010101010101;
12'd3436 : tab = 23'b10100011001110110000110;
12'd3437 : tab = 23'b10100011001010110111000;
12'd3438 : tab = 23'b10100011000110111101011;
12'd3439 : tab = 23'b10100011000011000011101;
12'd3440 : tab = 23'b10100010111111001010010;
12'd3441 : tab = 23'b10100010111011010000111;
12'd3442 : tab = 23'b10100010110111010111100;
12'd3443 : tab = 23'b10100010110011011110100;
12'd3444 : tab = 23'b10100010101111100101100;
12'd3445 : tab = 23'b10100010101011101100100;
12'd3446 : tab = 23'b10100010100111110011111;
12'd3447 : tab = 23'b10100010100011111011000;
12'd3448 : tab = 23'b10100010100000000010101;
12'd3449 : tab = 23'b10100010011100001010000;
12'd3450 : tab = 23'b10100010011000010001110;
12'd3451 : tab = 23'b10100010010100011001100;
12'd3452 : tab = 23'b10100010010000100001010;
12'd3453 : tab = 23'b10100010001100101001000;
12'd3454 : tab = 23'b10100010001000110001001;
12'd3455 : tab = 23'b10100010000100111001010;
12'd3456 : tab = 23'b10100010000001000001110;
12'd3457 : tab = 23'b10100001111101001010000;
12'd3458 : tab = 23'b10100001111001010010100;
12'd3459 : tab = 23'b10100001110101011011010;
12'd3460 : tab = 23'b10100001110001100011110;
12'd3461 : tab = 23'b10100001101101101100101;
12'd3462 : tab = 23'b10100001101001110101100;
12'd3463 : tab = 23'b10100001100101111110011;
12'd3464 : tab = 23'b10100001100010000111101;
12'd3465 : tab = 23'b10100001011110010000111;
12'd3466 : tab = 23'b10100001011010011010001;
12'd3467 : tab = 23'b10100001010110100011110;
12'd3468 : tab = 23'b10100001010010101101010;
12'd3469 : tab = 23'b10100001001110110111000;
12'd3470 : tab = 23'b10100001001011000000101;
12'd3471 : tab = 23'b10100001000111001010101;
12'd3472 : tab = 23'b10100001000011010100100;
12'd3473 : tab = 23'b10100000111111011110101;
12'd3474 : tab = 23'b10100000111011101000110;
12'd3475 : tab = 23'b10100000110111110011000;
12'd3476 : tab = 23'b10100000110011111101011;
12'd3477 : tab = 23'b10100000110000001000001;
12'd3478 : tab = 23'b10100000101100010010100;
12'd3479 : tab = 23'b10100000101000011101010;
12'd3480 : tab = 23'b10100000100100101000010;
12'd3481 : tab = 23'b10100000100000110011001;
12'd3482 : tab = 23'b10100000011100111110000;
12'd3483 : tab = 23'b10100000011001001001011;
12'd3484 : tab = 23'b10100000010101010100100;
12'd3485 : tab = 23'b10100000010001011111110;
12'd3486 : tab = 23'b10100000001101101011010;
12'd3487 : tab = 23'b10100000001001110111000;
12'd3488 : tab = 23'b10100000000110000010100;
12'd3489 : tab = 23'b10100000000010001110011;
12'd3490 : tab = 23'b10011111111110011010010;
12'd3491 : tab = 23'b10011111111010100110001;
12'd3492 : tab = 23'b10011111110110110010011;
12'd3493 : tab = 23'b10011111110010111110100;
12'd3494 : tab = 23'b10011111101111001010111;
12'd3495 : tab = 23'b10011111101011010111001;
12'd3496 : tab = 23'b10011111100111100011110;
12'd3497 : tab = 23'b10011111100011110000011;
12'd3498 : tab = 23'b10011111011111111101000;
12'd3499 : tab = 23'b10011111011100001001110;
12'd3500 : tab = 23'b10011111011000010110110;
12'd3501 : tab = 23'b10011111010100100011101;
12'd3502 : tab = 23'b10011111010000110001000;
12'd3503 : tab = 23'b10011111001100111110010;
12'd3504 : tab = 23'b10011111001001001011011;
12'd3505 : tab = 23'b10011111000101011001001;
12'd3506 : tab = 23'b10011111000001100110100;
12'd3507 : tab = 23'b10011110111101110100010;
12'd3508 : tab = 23'b10011110111010000010000;
12'd3509 : tab = 23'b10011110110110001111110;
12'd3510 : tab = 23'b10011110110010011101110;
12'd3511 : tab = 23'b10011110101110101011110;
12'd3512 : tab = 23'b10011110101010111010001;
12'd3513 : tab = 23'b10011110100111001000010;
12'd3514 : tab = 23'b10011110100011010110100;
12'd3515 : tab = 23'b10011110011111100101000;
12'd3516 : tab = 23'b10011110011011110011110;
12'd3517 : tab = 23'b10011110011000000010010;
12'd3518 : tab = 23'b10011110010100010001001;
12'd3519 : tab = 23'b10011110010000100000000;
12'd3520 : tab = 23'b10011110001100101111010;
12'd3521 : tab = 23'b10011110001000111110001;
12'd3522 : tab = 23'b10011110000101001101011;
12'd3523 : tab = 23'b10011110000001011100101;
12'd3524 : tab = 23'b10011101111101101100000;
12'd3525 : tab = 23'b10011101111001111011100;
12'd3526 : tab = 23'b10011101110110001011001;
12'd3527 : tab = 23'b10011101110010011010110;
12'd3528 : tab = 23'b10011101101110101010110;
12'd3529 : tab = 23'b10011101101010111010110;
12'd3530 : tab = 23'b10011101100111001010110;
12'd3531 : tab = 23'b10011101100011011010110;
12'd3532 : tab = 23'b10011101011111101011000;
12'd3533 : tab = 23'b10011101011011111011010;
12'd3534 : tab = 23'b10011101011000001011111;
12'd3535 : tab = 23'b10011101010100011100010;
12'd3536 : tab = 23'b10011101010000101101000;
12'd3537 : tab = 23'b10011101001100111101110;
12'd3538 : tab = 23'b10011101001001001110100;
12'd3539 : tab = 23'b10011101000101011111010;
12'd3540 : tab = 23'b10011101000001110000011;
12'd3541 : tab = 23'b10011100111110000001100;
12'd3542 : tab = 23'b10011100111010010010110;
12'd3543 : tab = 23'b10011100110110100100001;
12'd3544 : tab = 23'b10011100110010110101101;
12'd3545 : tab = 23'b10011100101111000111001;
12'd3546 : tab = 23'b10011100101011011000101;
12'd3547 : tab = 23'b10011100100111101010100;
12'd3548 : tab = 23'b10011100100011111100011;
12'd3549 : tab = 23'b10011100100000001110010;
12'd3550 : tab = 23'b10011100011100100000001;
12'd3551 : tab = 23'b10011100011000110010011;
12'd3552 : tab = 23'b10011100010101000100101;
12'd3553 : tab = 23'b10011100010001010110111;
12'd3554 : tab = 23'b10011100001101101001100;
12'd3555 : tab = 23'b10011100001001111100001;
12'd3556 : tab = 23'b10011100000110001110110;
12'd3557 : tab = 23'b10011100000010100001011;
12'd3558 : tab = 23'b10011011111110110100011;
12'd3559 : tab = 23'b10011011111011000111010;
12'd3560 : tab = 23'b10011011110111011010011;
12'd3561 : tab = 23'b10011011110011101101011;
12'd3562 : tab = 23'b10011011110000000000100;
12'd3563 : tab = 23'b10011011101100010100000;
12'd3564 : tab = 23'b10011011101000100111100;
12'd3565 : tab = 23'b10011011100100111010111;
12'd3566 : tab = 23'b10011011100001001110101;
12'd3567 : tab = 23'b10011011011101100010011;
12'd3568 : tab = 23'b10011011011001110110001;
12'd3569 : tab = 23'b10011011010110001010010;
12'd3570 : tab = 23'b10011011010010011110010;
12'd3571 : tab = 23'b10011011001110110010010;
12'd3572 : tab = 23'b10011011001011000110101;
12'd3573 : tab = 23'b10011011000111011010110;
12'd3574 : tab = 23'b10011011000011101111010;
12'd3575 : tab = 23'b10011011000000000011110;
12'd3576 : tab = 23'b10011010111100011000100;
12'd3577 : tab = 23'b10011010111000101101001;
12'd3578 : tab = 23'b10011010110101000010000;
12'd3579 : tab = 23'b10011010110001010110111;
12'd3580 : tab = 23'b10011010101101101100001;
12'd3581 : tab = 23'b10011010101010000001000;
12'd3582 : tab = 23'b10011010100110010110010;
12'd3583 : tab = 23'b10011010100010101011110;
12'd3584 : tab = 23'b10011010011111000001001;
12'd3585 : tab = 23'b10011010011011010110100;
12'd3586 : tab = 23'b10011010010111101100010;
12'd3587 : tab = 23'b10011010010100000010000;
12'd3588 : tab = 23'b10011010010000010111110;
12'd3589 : tab = 23'b10011010001100101101101;
12'd3590 : tab = 23'b10011010001001000011101;
12'd3591 : tab = 23'b10011010000101011001110;
12'd3592 : tab = 23'b10011010000001110000000;
12'd3593 : tab = 23'b10011001111110000110011;
12'd3594 : tab = 23'b10011001111010011100110;
12'd3595 : tab = 23'b10011001110110110011001;
12'd3596 : tab = 23'b10011001110011001001111;
12'd3597 : tab = 23'b10011001101111100000100;
12'd3598 : tab = 23'b10011001101011110111011;
12'd3599 : tab = 23'b10011001101000001110001;
12'd3600 : tab = 23'b10011001100100100101010;
12'd3601 : tab = 23'b10011001100000111100010;
12'd3602 : tab = 23'b10011001011101010011100;
12'd3603 : tab = 23'b10011001011001101010101;
12'd3604 : tab = 23'b10011001010110000010001;
12'd3605 : tab = 23'b10011001010010011001101;
12'd3606 : tab = 23'b10011001001110110001001;
12'd3607 : tab = 23'b10011001001011001000101;
12'd3608 : tab = 23'b10011001000111100000100;
12'd3609 : tab = 23'b10011001000011111000011;
12'd3610 : tab = 23'b10011001000000010000010;
12'd3611 : tab = 23'b10011000111100101000010;
12'd3612 : tab = 23'b10011000111001000000011;
12'd3613 : tab = 23'b10011000110101011000110;
12'd3614 : tab = 23'b10011000110001110001000;
12'd3615 : tab = 23'b10011000101110001001100;
12'd3616 : tab = 23'b10011000101010100010000;
12'd3617 : tab = 23'b10011000100110111010110;
12'd3618 : tab = 23'b10011000100011010011011;
12'd3619 : tab = 23'b10011000011111101100010;
12'd3620 : tab = 23'b10011000011100000101010;
12'd3621 : tab = 23'b10011000011000011110010;
12'd3622 : tab = 23'b10011000010100110111010;
12'd3623 : tab = 23'b10011000010001010000011;
12'd3624 : tab = 23'b10011000001101101001110;
12'd3625 : tab = 23'b10011000001010000011001;
12'd3626 : tab = 23'b10011000000110011100100;
12'd3627 : tab = 23'b10011000000010110110010;
12'd3628 : tab = 23'b10010111111111001111110;
12'd3629 : tab = 23'b10010111111011101001100;
12'd3630 : tab = 23'b10010111111000000011100;
12'd3631 : tab = 23'b10010111110100011101100;
12'd3632 : tab = 23'b10010111110000110111011;
12'd3633 : tab = 23'b10010111101101010001100;
12'd3634 : tab = 23'b10010111101001101100000;
12'd3635 : tab = 23'b10010111100110000110001;
12'd3636 : tab = 23'b10010111100010100000101;
12'd3637 : tab = 23'b10010111011110111011001;
12'd3638 : tab = 23'b10010111011011010101110;
12'd3639 : tab = 23'b10010111010111110000100;
12'd3640 : tab = 23'b10010111010100001011011;
12'd3641 : tab = 23'b10010111010000100110010;
12'd3642 : tab = 23'b10010111001101000001001;
12'd3643 : tab = 23'b10010111001001011100011;
12'd3644 : tab = 23'b10010111000101110111101;
12'd3645 : tab = 23'b10010111000010010010111;
12'd3646 : tab = 23'b10010110111110101110001;
12'd3647 : tab = 23'b10010110111011001001110;
12'd3648 : tab = 23'b10010110110111100101010;
12'd3649 : tab = 23'b10010110110100000001000;
12'd3650 : tab = 23'b10010110110000011100101;
12'd3651 : tab = 23'b10010110101100111000101;
12'd3652 : tab = 23'b10010110101001010100100;
12'd3653 : tab = 23'b10010110100101110000101;
12'd3654 : tab = 23'b10010110100010001100101;
12'd3655 : tab = 23'b10010110011110101000110;
12'd3656 : tab = 23'b10010110011011000101010;
12'd3657 : tab = 23'b10010110010111100001100;
12'd3658 : tab = 23'b10010110010011111110001;
12'd3659 : tab = 23'b10010110010000011010110;
12'd3660 : tab = 23'b10010110001100110111100;
12'd3661 : tab = 23'b10010110001001010100000;
12'd3662 : tab = 23'b10010110000101110001001;
12'd3663 : tab = 23'b10010110000010001101111;
12'd3664 : tab = 23'b10010101111110101011000;
12'd3665 : tab = 23'b10010101111011001000001;
12'd3666 : tab = 23'b10010101110111100101101;
12'd3667 : tab = 23'b10010101110100000010110;
12'd3668 : tab = 23'b10010101110000100000010;
12'd3669 : tab = 23'b10010101101100111101110;
12'd3670 : tab = 23'b10010101101001011011010;
12'd3671 : tab = 23'b10010101100101111001001;
12'd3672 : tab = 23'b10010101100010010110110;
12'd3673 : tab = 23'b10010101011110110100111;
12'd3674 : tab = 23'b10010101011011010010110;
12'd3675 : tab = 23'b10010101010111110001000;
12'd3676 : tab = 23'b10010101010100001111000;
12'd3677 : tab = 23'b10010101010000101101010;
12'd3678 : tab = 23'b10010101001101001011110;
12'd3679 : tab = 23'b10010101001001101010000;
12'd3680 : tab = 23'b10010101000110001000101;
12'd3681 : tab = 23'b10010101000010100111010;
12'd3682 : tab = 23'b10010100111111000101111;
12'd3683 : tab = 23'b10010100111011100100111;
12'd3684 : tab = 23'b10010100111000000011110;
12'd3685 : tab = 23'b10010100110100100010110;
12'd3686 : tab = 23'b10010100110001000001111;
12'd3687 : tab = 23'b10010100101101100000111;
12'd3688 : tab = 23'b10010100101010000000010;
12'd3689 : tab = 23'b10010100100110011111101;
12'd3690 : tab = 23'b10010100100010111111000;
12'd3691 : tab = 23'b10010100011111011110100;
12'd3692 : tab = 23'b10010100011011111110001;
12'd3693 : tab = 23'b10010100011000011101111;
12'd3694 : tab = 23'b10010100010100111101101;
12'd3695 : tab = 23'b10010100010001011101110;
12'd3696 : tab = 23'b10010100001101111101110;
12'd3697 : tab = 23'b10010100001010011101110;
12'd3698 : tab = 23'b10010100000110111110000;
12'd3699 : tab = 23'b10010100000011011110010;
12'd3700 : tab = 23'b10010011111111111110100;
12'd3701 : tab = 23'b10010011111100011111000;
12'd3702 : tab = 23'b10010011111000111111110;
12'd3703 : tab = 23'b10010011110101100000010;
12'd3704 : tab = 23'b10010011110010000001000;
12'd3705 : tab = 23'b10010011101110100001110;
12'd3706 : tab = 23'b10010011101011000010111;
12'd3707 : tab = 23'b10010011100111100011110;
12'd3708 : tab = 23'b10010011100100000100110;
12'd3709 : tab = 23'b10010011100000100101111;
12'd3710 : tab = 23'b10010011011101000111001;
12'd3711 : tab = 23'b10010011011001101000110;
12'd3712 : tab = 23'b10010011010110001010000;
12'd3713 : tab = 23'b10010011010010101011101;
12'd3714 : tab = 23'b10010011001111001101010;
12'd3715 : tab = 23'b10010011001011101110111;
12'd3716 : tab = 23'b10010011001000010000111;
12'd3717 : tab = 23'b10010011000100110010110;
12'd3718 : tab = 23'b10010011000001010100100;
12'd3719 : tab = 23'b10010010111101110110110;
12'd3720 : tab = 23'b10010010111010011000111;
12'd3721 : tab = 23'b10010010110110111011000;
12'd3722 : tab = 23'b10010010110011011101101;
12'd3723 : tab = 23'b10010010110000000000000;
12'd3724 : tab = 23'b10010010101100100010011;
12'd3725 : tab = 23'b10010010101001000101001;
12'd3726 : tab = 23'b10010010100101100111110;
12'd3727 : tab = 23'b10010010100010001010101;
12'd3728 : tab = 23'b10010010011110101101011;
12'd3729 : tab = 23'b10010010011011010000100;
12'd3730 : tab = 23'b10010010010111110011100;
12'd3731 : tab = 23'b10010010010100010110110;
12'd3732 : tab = 23'b10010010010000111001111;
12'd3733 : tab = 23'b10010010001101011101010;
12'd3734 : tab = 23'b10010010001010000000100;
12'd3735 : tab = 23'b10010010000110100100000;
12'd3736 : tab = 23'b10010010000011000111111;
12'd3737 : tab = 23'b10010001111111101011011;
12'd3738 : tab = 23'b10010001111100001111000;
12'd3739 : tab = 23'b10010001111000110011001;
12'd3740 : tab = 23'b10010001110101010111000;
12'd3741 : tab = 23'b10010001110001111010111;
12'd3742 : tab = 23'b10010001101110011111001;
12'd3743 : tab = 23'b10010001101011000011011;
12'd3744 : tab = 23'b10010001100111100111101;
12'd3745 : tab = 23'b10010001100100001011111;
12'd3746 : tab = 23'b10010001100000110000100;
12'd3747 : tab = 23'b10010001011101010101000;
12'd3748 : tab = 23'b10010001011001111001110;
12'd3749 : tab = 23'b10010001010110011110011;
12'd3750 : tab = 23'b10010001010011000011010;
12'd3751 : tab = 23'b10010001001111101000000;
12'd3752 : tab = 23'b10010001001100001101000;
12'd3753 : tab = 23'b10010001001000110010000;
12'd3754 : tab = 23'b10010001000101010111011;
12'd3755 : tab = 23'b10010001000001111100110;
12'd3756 : tab = 23'b10010000111110100010001;
12'd3757 : tab = 23'b10010000111011000111100;
12'd3758 : tab = 23'b10010000110111101100111;
12'd3759 : tab = 23'b10010000110100010010101;
12'd3760 : tab = 23'b10010000110000111000010;
12'd3761 : tab = 23'b10010000101101011110001;
12'd3762 : tab = 23'b10010000101010000011111;
12'd3763 : tab = 23'b10010000100110101001110;
12'd3764 : tab = 23'b10010000100011010000000;
12'd3765 : tab = 23'b10010000011111110110000;
12'd3766 : tab = 23'b10010000011100011100011;
12'd3767 : tab = 23'b10010000011001000010100;
12'd3768 : tab = 23'b10010000010101101001000;
12'd3769 : tab = 23'b10010000010010001111100;
12'd3770 : tab = 23'b10010000001110110110000;
12'd3771 : tab = 23'b10010000001011011100110;
12'd3772 : tab = 23'b10010000001000000011011;
12'd3773 : tab = 23'b10010000000100101010010;
12'd3774 : tab = 23'b10010000000001010001001;
12'd3775 : tab = 23'b10001111111101111000000;
12'd3776 : tab = 23'b10001111111010011111010;
12'd3777 : tab = 23'b10001111110111000110010;
12'd3778 : tab = 23'b10001111110011101101110;
12'd3779 : tab = 23'b10001111110000010101000;
12'd3780 : tab = 23'b10001111101100111100100;
12'd3781 : tab = 23'b10001111101001100011111;
12'd3782 : tab = 23'b10001111100110001011100;
12'd3783 : tab = 23'b10001111100010110011001;
12'd3784 : tab = 23'b10001111011111011011001;
12'd3785 : tab = 23'b10001111011100000010110;
12'd3786 : tab = 23'b10001111011000101010110;
12'd3787 : tab = 23'b10001111010101010010110;
12'd3788 : tab = 23'b10001111010001111010110;
12'd3789 : tab = 23'b10001111001110100011001;
12'd3790 : tab = 23'b10001111001011001011010;
12'd3791 : tab = 23'b10001111000111110011110;
12'd3792 : tab = 23'b10001111000100011100010;
12'd3793 : tab = 23'b10001111000001000100101;
12'd3794 : tab = 23'b10001110111101101101011;
12'd3795 : tab = 23'b10001110111010010110001;
12'd3796 : tab = 23'b10001110110110111110111;
12'd3797 : tab = 23'b10001110110011100111101;
12'd3798 : tab = 23'b10001110110000010000110;
12'd3799 : tab = 23'b10001110101100111001110;
12'd3800 : tab = 23'b10001110101001100011000;
12'd3801 : tab = 23'b10001110100110001100001;
12'd3802 : tab = 23'b10001110100010110101100;
12'd3803 : tab = 23'b10001110011111011110110;
12'd3804 : tab = 23'b10001110011100001000010;
12'd3805 : tab = 23'b10001110011000110001110;
12'd3806 : tab = 23'b10001110010101011011101;
12'd3807 : tab = 23'b10001110010010000101001;
12'd3808 : tab = 23'b10001110001110101111000;
12'd3809 : tab = 23'b10001110001011011000111;
12'd3810 : tab = 23'b10001110001000000010110;
12'd3811 : tab = 23'b10001110000100101101000;
12'd3812 : tab = 23'b10001110000001010111000;
12'd3813 : tab = 23'b10001101111110000001100;
12'd3814 : tab = 23'b10001101111010101011110;
12'd3815 : tab = 23'b10001101110111010110000;
12'd3816 : tab = 23'b10001101110100000000101;
12'd3817 : tab = 23'b10001101110000101011000;
12'd3818 : tab = 23'b10001101101101010101111;
12'd3819 : tab = 23'b10001101101010000000100;
12'd3820 : tab = 23'b10001101100110101011010;
12'd3821 : tab = 23'b10001101100011010110001;
12'd3822 : tab = 23'b10001101100000000001001;
12'd3823 : tab = 23'b10001101011100101100001;
12'd3824 : tab = 23'b10001101011001010111100;
12'd3825 : tab = 23'b10001101010110000010110;
12'd3826 : tab = 23'b10001101010010101110000;
12'd3827 : tab = 23'b10001101001111011001100;
12'd3828 : tab = 23'b10001101001100000101000;
12'd3829 : tab = 23'b10001101001000110000011;
12'd3830 : tab = 23'b10001101000101011100001;
12'd3831 : tab = 23'b10001101000010000111111;
12'd3832 : tab = 23'b10001100111110110011101;
12'd3833 : tab = 23'b10001100111011011111100;
12'd3834 : tab = 23'b10001100111000001011100;
12'd3835 : tab = 23'b10001100110100110111101;
12'd3836 : tab = 23'b10001100110001100011110;
12'd3837 : tab = 23'b10001100101110001111111;
12'd3838 : tab = 23'b10001100101010111100011;
12'd3839 : tab = 23'b10001100100111101000111;
12'd3840 : tab = 23'b10001100100100010101011;
12'd3841 : tab = 23'b10001100100001000001111;
12'd3842 : tab = 23'b10001100011101101110011;
12'd3843 : tab = 23'b10001100011010011011010;
12'd3844 : tab = 23'b10001100010111001000001;
12'd3845 : tab = 23'b10001100010011110101000;
12'd3846 : tab = 23'b10001100010000100001111;
12'd3847 : tab = 23'b10001100001101001110110;
12'd3848 : tab = 23'b10001100001001111100000;
12'd3849 : tab = 23'b10001100000110101001010;
12'd3850 : tab = 23'b10001100000011010110100;
12'd3851 : tab = 23'b10001100000000000100001;
12'd3852 : tab = 23'b10001011111100110001011;
12'd3853 : tab = 23'b10001011111001011111000;
12'd3854 : tab = 23'b10001011110110001100101;
12'd3855 : tab = 23'b10001011110010111010010;
12'd3856 : tab = 23'b10001011101111101000010;
12'd3857 : tab = 23'b10001011101100010110000;
12'd3858 : tab = 23'b10001011101001000100000;
12'd3859 : tab = 23'b10001011100101110010010;
12'd3860 : tab = 23'b10001011100010100000010;
12'd3861 : tab = 23'b10001011011111001110100;
12'd3862 : tab = 23'b10001011011011111100101;
12'd3863 : tab = 23'b10001011011000101011000;
12'd3864 : tab = 23'b10001011010101011001011;
12'd3865 : tab = 23'b10001011010010001000001;
12'd3866 : tab = 23'b10001011001110110110110;
12'd3867 : tab = 23'b10001011001011100101010;
12'd3868 : tab = 23'b10001011001000010100000;
12'd3869 : tab = 23'b10001011000101000011000;
12'd3870 : tab = 23'b10001011000001110001111;
12'd3871 : tab = 23'b10001010111110100001000;
12'd3872 : tab = 23'b10001010111011010000001;
12'd3873 : tab = 23'b10001010110111111111010;
12'd3874 : tab = 23'b10001010110100101110011;
12'd3875 : tab = 23'b10001010110001011101111;
12'd3876 : tab = 23'b10001010101110001101010;
12'd3877 : tab = 23'b10001010101010111100111;
12'd3878 : tab = 23'b10001010100111101100011;
12'd3879 : tab = 23'b10001010100100011100000;
12'd3880 : tab = 23'b10001010100001001011110;
12'd3881 : tab = 23'b10001010011101111011101;
12'd3882 : tab = 23'b10001010011010101011100;
12'd3883 : tab = 23'b10001010010111011011011;
12'd3884 : tab = 23'b10001010010100001011101;
12'd3885 : tab = 23'b10001010010000111011110;
12'd3886 : tab = 23'b10001010001101101100000;
12'd3887 : tab = 23'b10001010001010011100010;
12'd3888 : tab = 23'b10001010000111001100101;
12'd3889 : tab = 23'b10001010000011111101000;
12'd3890 : tab = 23'b10001010000000101101100;
12'd3891 : tab = 23'b10001001111101011110001;
12'd3892 : tab = 23'b10001001111010001111000;
12'd3893 : tab = 23'b10001001110110111111110;
12'd3894 : tab = 23'b10001001110011110000100;
12'd3895 : tab = 23'b10001001110000100001100;
12'd3896 : tab = 23'b10001001101101010010110;
12'd3897 : tab = 23'b10001001101010000011110;
12'd3898 : tab = 23'b10001001100110110100110;
12'd3899 : tab = 23'b10001001100011100110001;
12'd3900 : tab = 23'b10001001100000010111100;
12'd3901 : tab = 23'b10001001011101001000111;
12'd3902 : tab = 23'b10001001011001111010100;
12'd3903 : tab = 23'b10001001010110101100000;
12'd3904 : tab = 23'b10001001010011011101100;
12'd3905 : tab = 23'b10001001010000001111100;
12'd3906 : tab = 23'b10001001001101000001010;
12'd3907 : tab = 23'b10001001001001110011000;
12'd3908 : tab = 23'b10001001000110100101001;
12'd3909 : tab = 23'b10001001000011010111010;
12'd3910 : tab = 23'b10001001000000001001011;
12'd3911 : tab = 23'b10001000111100111011100;
12'd3912 : tab = 23'b10001000111001101101110;
12'd3913 : tab = 23'b10001000110110100000001;
12'd3914 : tab = 23'b10001000110011010010101;
12'd3915 : tab = 23'b10001000110000000101001;
12'd3916 : tab = 23'b10001000101100111000000;
12'd3917 : tab = 23'b10001000101001101010100;
12'd3918 : tab = 23'b10001000100110011101011;
12'd3919 : tab = 23'b10001000100011010000000;
12'd3920 : tab = 23'b10001000100000000011001;
12'd3921 : tab = 23'b10001000011100110110000;
12'd3922 : tab = 23'b10001000011001101001000;
12'd3923 : tab = 23'b10001000010110011100010;
12'd3924 : tab = 23'b10001000010011001111100;
12'd3925 : tab = 23'b10001000010000000010110;
12'd3926 : tab = 23'b10001000001100110110010;
12'd3927 : tab = 23'b10001000001001101001110;
12'd3928 : tab = 23'b10001000000110011101001;
12'd3929 : tab = 23'b10001000000011010000110;
12'd3930 : tab = 23'b10001000000000000100110;
12'd3931 : tab = 23'b10000111111100111000011;
12'd3932 : tab = 23'b10000111111001101100010;
12'd3933 : tab = 23'b10000111110110100000010;
12'd3934 : tab = 23'b10000111110011010100010;
12'd3935 : tab = 23'b10000111110000001000011;
12'd3936 : tab = 23'b10000111101100111100011;
12'd3937 : tab = 23'b10000111101001110000110;
12'd3938 : tab = 23'b10000111100110100101001;
12'd3939 : tab = 23'b10000111100011011001100;
12'd3940 : tab = 23'b10000111100000001101111;
12'd3941 : tab = 23'b10000111011101000010100;
12'd3942 : tab = 23'b10000111011001110111010;
12'd3943 : tab = 23'b10000111010110101011110;
12'd3944 : tab = 23'b10000111010011100000110;
12'd3945 : tab = 23'b10000111010000010101101;
12'd3946 : tab = 23'b10000111001101001010011;
12'd3947 : tab = 23'b10000111001001111111100;
12'd3948 : tab = 23'b10000111000110110100101;
12'd3949 : tab = 23'b10000111000011101001110;
12'd3950 : tab = 23'b10000111000000011110111;
12'd3951 : tab = 23'b10000110111101010100011;
12'd3952 : tab = 23'b10000110111010001001111;
12'd3953 : tab = 23'b10000110110110111111011;
12'd3954 : tab = 23'b10000110110011110100111;
12'd3955 : tab = 23'b10000110110000101010011;
12'd3956 : tab = 23'b10000110101101100000010;
12'd3957 : tab = 23'b10000110101010010110000;
12'd3958 : tab = 23'b10000110100111001100000;
12'd3959 : tab = 23'b10000110100100000001111;
12'd3960 : tab = 23'b10000110100000110111110;
12'd3961 : tab = 23'b10000110011101101110000;
12'd3962 : tab = 23'b10000110011010100100000;
12'd3963 : tab = 23'b10000110010111011010010;
12'd3964 : tab = 23'b10000110010100010000110;
12'd3965 : tab = 23'b10000110010001000111000;
12'd3966 : tab = 23'b10000110001101111101101;
12'd3967 : tab = 23'b10000110001010110100010;
12'd3968 : tab = 23'b10000110000111101010111;
12'd3969 : tab = 23'b10000110000100100001100;
12'd3970 : tab = 23'b10000110000001011000001;
12'd3971 : tab = 23'b10000101111110001111001;
12'd3972 : tab = 23'b10000101111011000110001;
12'd3973 : tab = 23'b10000101110111111101001;
12'd3974 : tab = 23'b10000101110100110100001;
12'd3975 : tab = 23'b10000101110001101011100;
12'd3976 : tab = 23'b10000101101110100010110;
12'd3977 : tab = 23'b10000101101011011001111;
12'd3978 : tab = 23'b10000101101000010001010;
12'd3979 : tab = 23'b10000101100101001000101;
12'd3980 : tab = 23'b10000101100010000000011;
12'd3981 : tab = 23'b10000101011110111000000;
12'd3982 : tab = 23'b10000101011011101111110;
12'd3983 : tab = 23'b10000101011000100111100;
12'd3984 : tab = 23'b10000101010101011111011;
12'd3985 : tab = 23'b10000101010010010111001;
12'd3986 : tab = 23'b10000101001111001111010;
12'd3987 : tab = 23'b10000101001100000111010;
12'd3988 : tab = 23'b10000101001000111111100;
12'd3989 : tab = 23'b10000101000101110111101;
12'd3990 : tab = 23'b10000101000010110000000;
12'd3991 : tab = 23'b10000100111111101000010;
12'd3992 : tab = 23'b10000100111100100000110;
12'd3993 : tab = 23'b10000100111001011001010;
12'd3994 : tab = 23'b10000100110110010001110;
12'd3995 : tab = 23'b10000100110011001010101;
12'd3996 : tab = 23'b10000100110000000011010;
12'd3997 : tab = 23'b10000100101100111100000;
12'd3998 : tab = 23'b10000100101001110100111;
12'd3999 : tab = 23'b10000100100110101110001;
12'd4000 : tab = 23'b10000100100011100111000;
12'd4001 : tab = 23'b10000100100000100000000;
12'd4002 : tab = 23'b10000100011101011001010;
12'd4003 : tab = 23'b10000100011010010010110;
12'd4004 : tab = 23'b10000100010111001100000;
12'd4005 : tab = 23'b10000100010100000101010;
12'd4006 : tab = 23'b10000100010000111110111;
12'd4007 : tab = 23'b10000100001101111000100;
12'd4008 : tab = 23'b10000100001010110010001;
12'd4009 : tab = 23'b10000100000111101011110;
12'd4010 : tab = 23'b10000100000100100101100;
12'd4011 : tab = 23'b10000100000001011111011;
12'd4012 : tab = 23'b10000011111110011001011;
12'd4013 : tab = 23'b10000011111011010011011;
12'd4014 : tab = 23'b10000011111000001101011;
12'd4015 : tab = 23'b10000011110101000111110;
12'd4016 : tab = 23'b10000011110010000001110;
12'd4017 : tab = 23'b10000011101110111100001;
12'd4018 : tab = 23'b10000011101011110110100;
12'd4019 : tab = 23'b10000011101000110000111;
12'd4020 : tab = 23'b10000011100101101011101;
12'd4021 : tab = 23'b10000011100010100110010;
12'd4022 : tab = 23'b10000011011111100001000;
12'd4023 : tab = 23'b10000011011100011011100;
12'd4024 : tab = 23'b10000011011001010110100;
12'd4025 : tab = 23'b10000011010110010001011;
12'd4026 : tab = 23'b10000011010011001100010;
12'd4027 : tab = 23'b10000011010000000111010;
12'd4028 : tab = 23'b10000011001101000010011;
12'd4029 : tab = 23'b10000011001001111101100;
12'd4030 : tab = 23'b10000011000110111001000;
12'd4031 : tab = 23'b10000011000011110100010;
12'd4032 : tab = 23'b10000011000000101111101;
12'd4033 : tab = 23'b10000010111101101011001;
12'd4034 : tab = 23'b10000010111010100110101;
12'd4035 : tab = 23'b10000010110111100010100;
12'd4036 : tab = 23'b10000010110100011110000;
12'd4037 : tab = 23'b10000010110001011001111;
12'd4038 : tab = 23'b10000010101110010101110;
12'd4039 : tab = 23'b10000010101011010001101;
12'd4040 : tab = 23'b10000010101000001101100;
12'd4041 : tab = 23'b10000010100101001001110;
12'd4042 : tab = 23'b10000010100010000101110;
12'd4043 : tab = 23'b10000010011111000001111;
12'd4044 : tab = 23'b10000010011011111110001;
12'd4045 : tab = 23'b10000010011000111010110;
12'd4046 : tab = 23'b10000010010101110111000;
12'd4047 : tab = 23'b10000010010010110011101;
12'd4048 : tab = 23'b10000010001111110000000;
12'd4049 : tab = 23'b10000010001100101100111;
12'd4050 : tab = 23'b10000010001001101001100;
12'd4051 : tab = 23'b10000010000110100110010;
12'd4052 : tab = 23'b10000010000011100011001;
12'd4053 : tab = 23'b10000010000000100000001;
12'd4054 : tab = 23'b10000001111101011101001;
12'd4055 : tab = 23'b10000001111010011010001;
12'd4056 : tab = 23'b10000001110111010111010;
12'd4057 : tab = 23'b10000001110100010100100;
12'd4058 : tab = 23'b10000001110001010001111;
12'd4059 : tab = 23'b10000001101110001111010;
12'd4060 : tab = 23'b10000001101011001100101;
12'd4061 : tab = 23'b10000001101000001010010;
12'd4062 : tab = 23'b10000001100101000111110;
12'd4063 : tab = 23'b10000001100010000101100;
12'd4064 : tab = 23'b10000001011111000011010;
12'd4065 : tab = 23'b10000001011100000001000;
12'd4066 : tab = 23'b10000001011000111110110;
12'd4067 : tab = 23'b10000001010101111100110;
12'd4068 : tab = 23'b10000001010010111010110;
12'd4069 : tab = 23'b10000001001111111000110;
12'd4070 : tab = 23'b10000001001100110111000;
12'd4071 : tab = 23'b10000001001001110101011;
12'd4072 : tab = 23'b10000001000110110011100;
12'd4073 : tab = 23'b10000001000011110001110;
12'd4074 : tab = 23'b10000001000000110000010;
12'd4075 : tab = 23'b10000000111101101111000;
12'd4076 : tab = 23'b10000000111010101101100;
12'd4077 : tab = 23'b10000000110111101100000;
12'd4078 : tab = 23'b10000000110100101010111;
12'd4079 : tab = 23'b10000000110001101001110;
12'd4080 : tab = 23'b10000000101110101000101;
12'd4081 : tab = 23'b10000000101011100111100;
12'd4082 : tab = 23'b10000000101000100110011;
12'd4083 : tab = 23'b10000000100101100101101;
12'd4084 : tab = 23'b10000000100010100100110;
12'd4085 : tab = 23'b10000000011111100100000;
12'd4086 : tab = 23'b10000000011100100011011;
12'd4087 : tab = 23'b10000000011001100010101;
12'd4088 : tab = 23'b10000000010110100010000;
12'd4089 : tab = 23'b10000000010011100001100;
12'd4090 : tab = 23'b10000000010000100001001;
12'd4091 : tab = 23'b10000000001101100000110;
12'd4092 : tab = 23'b10000000001010100000011;
12'd4093 : tab = 23'b10000000000111100000011;
12'd4094 : tab = 23'b10000000000100100000010;
12'd4095 : tab = 23'b10000000000001100000000;
  endcase
  end
  endfunction
  
  function [22:0] tab2 (
    input [11:0] N
  );
  begin
  case(N)
12'd0 : tab2 = 23'b11111111110100000000110;
12'd1 : tab2 = 23'b11111111011100000010010;
12'd2 : tab2 = 23'b11111111000100000110000;
12'd3 : tab2 = 23'b11111110101100001011010;
12'd4 : tab2 = 23'b11111110010100010011100;
12'd5 : tab2 = 23'b11111101111100011100100;
12'd6 : tab2 = 23'b11111101100100100111110;
12'd7 : tab2 = 23'b11111101001100110100100;
12'd8 : tab2 = 23'b11111100110101000100001;
12'd9 : tab2 = 23'b11111100011101010100101;
12'd10 : tab2 = 23'b11111100000101100111010;
12'd11 : tab2 = 23'b11111011101101111011011;
12'd12 : tab2 = 23'b11111011010110010001110;
12'd13 : tab2 = 23'b11111010111110101001100;
12'd14 : tab2 = 23'b11111010100111000100000;
12'd15 : tab2 = 23'b11111010001111011111010;
12'd16 : tab2 = 23'b11111001110111111101000;
12'd17 : tab2 = 23'b11111001100000011100100;
12'd18 : tab2 = 23'b11111001001000111101110;
12'd19 : tab2 = 23'b11111000110001100001000;
12'd20 : tab2 = 23'b11111000011010000101110;
12'd21 : tab2 = 23'b11111000000010101100110;
12'd22 : tab2 = 23'b11110111101011010100110;
12'd23 : tab2 = 23'b11110111010011111111100;
12'd24 : tab2 = 23'b11110110111100101011010;
12'd25 : tab2 = 23'b11110110100101011001001;
12'd26 : tab2 = 23'b11110110001110001001010;
12'd27 : tab2 = 23'b11110101110110111010001;
12'd28 : tab2 = 23'b11110101011111101101101;
12'd29 : tab2 = 23'b11110101001000100010110;
12'd30 : tab2 = 23'b11110100110001011001100;
12'd31 : tab2 = 23'b11110100011010010010000;
12'd32 : tab2 = 23'b11110100000011001100110;
12'd33 : tab2 = 23'b11110011101100001000111;
12'd34 : tab2 = 23'b11110011010101000110111;
12'd35 : tab2 = 23'b11110010111110000110101;
12'd36 : tab2 = 23'b11110010100111000111110;
12'd37 : tab2 = 23'b11110010010000001010111;
12'd38 : tab2 = 23'b11110001111001010000000;
12'd39 : tab2 = 23'b11110001100010010111001;
12'd40 : tab2 = 23'b11110001001011011111101;
12'd41 : tab2 = 23'b11110000110100101001100;
12'd42 : tab2 = 23'b11110000011101110101100;
12'd43 : tab2 = 23'b11110000000111000011000;
12'd44 : tab2 = 23'b11101111110000010010101;
12'd45 : tab2 = 23'b11101111011001100100001;
12'd46 : tab2 = 23'b11101111000010110110110;
12'd47 : tab2 = 23'b11101110101100001011110;
12'd48 : tab2 = 23'b11101110010101100010010;
12'd49 : tab2 = 23'b11101101111110111010100;
12'd50 : tab2 = 23'b11101101101000010100010;
12'd51 : tab2 = 23'b11101101010001110000000;
12'd52 : tab2 = 23'b11101100111011001101100;
12'd53 : tab2 = 23'b11101100100100101100000;
12'd54 : tab2 = 23'b11101100001110001101000;
12'd55 : tab2 = 23'b11101011110111101111011;
12'd56 : tab2 = 23'b11101011100001010011101;
12'd57 : tab2 = 23'b11101011001010111001101;
12'd58 : tab2 = 23'b11101010110100100000110;
12'd59 : tab2 = 23'b11101010011110001010011;
12'd60 : tab2 = 23'b11101010000111110101010;
12'd61 : tab2 = 23'b11101001110001100010001;
12'd62 : tab2 = 23'b11101001011011010000110;
12'd63 : tab2 = 23'b11101001000101000000011;
12'd64 : tab2 = 23'b11101000101110110010010;
12'd65 : tab2 = 23'b11101000011000100101110;
12'd66 : tab2 = 23'b11101000000010011010110;
12'd67 : tab2 = 23'b11100111101100010001100;
12'd68 : tab2 = 23'b11100111010110001001101;
12'd69 : tab2 = 23'b11100111000000000100010;
12'd70 : tab2 = 23'b11100110101001111111111;
12'd71 : tab2 = 23'b11100110010011111101010;
12'd72 : tab2 = 23'b11100101111101111100100;
12'd73 : tab2 = 23'b11100101100111111101001;
12'd74 : tab2 = 23'b11100101010001111111101;
12'd75 : tab2 = 23'b11100100111100000011011;
12'd76 : tab2 = 23'b11100100100110001001110;
12'd77 : tab2 = 23'b11100100010000010000101;
12'd78 : tab2 = 23'b11100011111010011001101;
12'd79 : tab2 = 23'b11100011100100100100101;
12'd80 : tab2 = 23'b11100011001110110000101;
12'd81 : tab2 = 23'b11100010111000111111001;
12'd82 : tab2 = 23'b11100010100011001110101;
12'd83 : tab2 = 23'b11100010001101011111100;
12'd84 : tab2 = 23'b11100001110111110010011;
12'd85 : tab2 = 23'b11100001100010000110110;
12'd86 : tab2 = 23'b11100001001100011101010;
12'd87 : tab2 = 23'b11100000110110110100110;
12'd88 : tab2 = 23'b11100000100001001101111;
12'd89 : tab2 = 23'b11100000001011101000110;
12'd90 : tab2 = 23'b11011111110110000101110;
12'd91 : tab2 = 23'b11011111100000100011011;
12'd92 : tab2 = 23'b11011111001011000011011;
12'd93 : tab2 = 23'b11011110110101100100110;
12'd94 : tab2 = 23'b11011110100000001000011;
12'd95 : tab2 = 23'b11011110001010101100011;
12'd96 : tab2 = 23'b11011101110101010011000;
12'd97 : tab2 = 23'b11011101011111111010100;
12'd98 : tab2 = 23'b11011101001010100011111;
12'd99 : tab2 = 23'b11011100110101001110111;
12'd100 : tab2 = 23'b11011100011111111011111;
12'd101 : tab2 = 23'b11011100001010101001101;
12'd102 : tab2 = 23'b11011011110101011001011;
12'd103 : tab2 = 23'b11011011100000001011001;
12'd104 : tab2 = 23'b11011011001010111101100;
12'd105 : tab2 = 23'b11011010110101110010001;
12'd106 : tab2 = 23'b11011010100000101000010;
12'd107 : tab2 = 23'b11011010001011011111110;
12'd108 : tab2 = 23'b11011001110110011001000;
12'd109 : tab2 = 23'b11011001100001010011111;
12'd110 : tab2 = 23'b11011001001100001111111;
12'd111 : tab2 = 23'b11011000110111001110001;
12'd112 : tab2 = 23'b11011000100010001101100;
12'd113 : tab2 = 23'b11011000001101001110001;
12'd114 : tab2 = 23'b11010111111000010000110;
12'd115 : tab2 = 23'b11010111100011010100110;
12'd116 : tab2 = 23'b11010111001110011010110;
12'd117 : tab2 = 23'b11010110111001100010001;
12'd118 : tab2 = 23'b11010110100100101010011;
12'd119 : tab2 = 23'b11010110001111110100110;
12'd120 : tab2 = 23'b11010101111011000000001;
12'd121 : tab2 = 23'b11010101100110001110010;
12'd122 : tab2 = 23'b11010101010001011100111;
12'd123 : tab2 = 23'b11010100111100101101010;
12'd124 : tab2 = 23'b11010100100111111111011;
12'd125 : tab2 = 23'b11010100010011010010011;
12'd126 : tab2 = 23'b11010011111110100111101;
12'd127 : tab2 = 23'b11010011101001111110011;
12'd128 : tab2 = 23'b11010011010101010110011;
12'd129 : tab2 = 23'b11010011000000101111101;
12'd130 : tab2 = 23'b11010010101100001011000;
12'd131 : tab2 = 23'b11010010010111100111010;
12'd132 : tab2 = 23'b11010010000011000101101;
12'd133 : tab2 = 23'b11010001101110100100110;
12'd134 : tab2 = 23'b11010001011010000110001;
12'd135 : tab2 = 23'b11010001000101101000110;
12'd136 : tab2 = 23'b11010000110001001100111;
12'd137 : tab2 = 23'b11010000011100110010011;
12'd138 : tab2 = 23'b11010000001000011000111;
12'd139 : tab2 = 23'b11001111110100000010001;
12'd140 : tab2 = 23'b11001111011111101011110;
12'd141 : tab2 = 23'b11001111001011010111010;
12'd142 : tab2 = 23'b11001110110111000100010;
12'd143 : tab2 = 23'b11001110100010110011000;
12'd144 : tab2 = 23'b11001110001110100010101;
12'd145 : tab2 = 23'b11001101111010010100010;
12'd146 : tab2 = 23'b11001101100110000111010;
12'd147 : tab2 = 23'b11001101010001111011110;
12'd148 : tab2 = 23'b11001100111101110001101;
12'd149 : tab2 = 23'b11001100101001101000011;
12'd150 : tab2 = 23'b11001100010101100001111;
12'd151 : tab2 = 23'b11001100000001011100000;
12'd152 : tab2 = 23'b11001011101101010111101;
12'd153 : tab2 = 23'b11001011011001010100101;
12'd154 : tab2 = 23'b11001011000101010011010;
12'd155 : tab2 = 23'b11001010110001010011001;
12'd156 : tab2 = 23'b11001010011101010101001;
12'd157 : tab2 = 23'b11001010001001011000001;
12'd158 : tab2 = 23'b11001001110101011100101;
12'd159 : tab2 = 23'b11001001100001100010001;
12'd160 : tab2 = 23'b11001001001101101001111;
12'd161 : tab2 = 23'b11001000111001110010001;
12'd162 : tab2 = 23'b11001000100101111100101;
12'd163 : tab2 = 23'b11001000010010001000001;
12'd164 : tab2 = 23'b11000111111110010101111;
12'd165 : tab2 = 23'b11000111101010100011111;
12'd166 : tab2 = 23'b11000111010110110011100;
12'd167 : tab2 = 23'b11000111000011000101001;
12'd168 : tab2 = 23'b11000110101111010111100;
12'd169 : tab2 = 23'b11000110011011101100000;
12'd170 : tab2 = 23'b11000110001000000001110;
12'd171 : tab2 = 23'b11000101110100011000101;
12'd172 : tab2 = 23'b11000101100000110000111;
12'd173 : tab2 = 23'b11000101001101001011000;
12'd174 : tab2 = 23'b11000100111001100110011;
12'd175 : tab2 = 23'b11000100100110000011001;
12'd176 : tab2 = 23'b11000100010010100001000;
12'd177 : tab2 = 23'b11000011111111000000100;
12'd178 : tab2 = 23'b11000011101011100001011;
12'd179 : tab2 = 23'b11000011011000000011110;
12'd180 : tab2 = 23'b11000011000100100111010;
12'd181 : tab2 = 23'b11000010110001001100100;
12'd182 : tab2 = 23'b11000010011101110011000;
12'd183 : tab2 = 23'b11000010001010011011001;
12'd184 : tab2 = 23'b11000001110111000100011;
12'd185 : tab2 = 23'b11000001100011101110111;
12'd186 : tab2 = 23'b11000001010000011010101;
12'd187 : tab2 = 23'b11000000111101001000010;
12'd188 : tab2 = 23'b11000000101001110111000;
12'd189 : tab2 = 23'b11000000010110100111100;
12'd190 : tab2 = 23'b11000000000011011000111;
12'd191 : tab2 = 23'b10111111110000001011100;
12'd192 : tab2 = 23'b10111111011101000000001;
12'd193 : tab2 = 23'b10111111001001110101111;
12'd194 : tab2 = 23'b10111110110110101100010;
12'd195 : tab2 = 23'b10111110100011100101001;
12'd196 : tab2 = 23'b10111110010000011110110;
12'd197 : tab2 = 23'b10111101111101011010001;
12'd198 : tab2 = 23'b10111101101010010110001;
12'd199 : tab2 = 23'b10111101010111010100000;
12'd200 : tab2 = 23'b10111101000100010011110;
12'd201 : tab2 = 23'b10111100110001010011101;
12'd202 : tab2 = 23'b10111100011110010101111;
12'd203 : tab2 = 23'b10111100001011011001000;
12'd204 : tab2 = 23'b10111011111000011101101;
12'd205 : tab2 = 23'b10111011100101100011010;
12'd206 : tab2 = 23'b10111011010010101010110;
12'd207 : tab2 = 23'b10111010111111110011101;
12'd208 : tab2 = 23'b10111010101100111101001;
12'd209 : tab2 = 23'b10111010011010001000101;
12'd210 : tab2 = 23'b10111010000111010101010;
12'd211 : tab2 = 23'b10111001110100100011001;
12'd212 : tab2 = 23'b10111001100001110010111;
12'd213 : tab2 = 23'b10111001001111000011001;
12'd214 : tab2 = 23'b10111000111100010100101;
12'd215 : tab2 = 23'b10111000101001101000000;
12'd216 : tab2 = 23'b10111000010110111100111;
12'd217 : tab2 = 23'b10111000000100010010011;
12'd218 : tab2 = 23'b10110111110001101010000;
12'd219 : tab2 = 23'b10110111011111000010010;
12'd220 : tab2 = 23'b10110111001100011100010;
12'd221 : tab2 = 23'b10110110111001110111100;
12'd222 : tab2 = 23'b10110110100111010100000;
12'd223 : tab2 = 23'b10110110010100110001101;
12'd224 : tab2 = 23'b10110110000010010000111;
12'd225 : tab2 = 23'b10110101101111110000101;
12'd226 : tab2 = 23'b10110101011101010010101;
12'd227 : tab2 = 23'b10110101001010110101110;
12'd228 : tab2 = 23'b10110100111000011001110;
12'd229 : tab2 = 23'b10110100100101111111100;
12'd230 : tab2 = 23'b10110100010011100110010;
12'd231 : tab2 = 23'b10110100000001001110001;
12'd232 : tab2 = 23'b10110011101110111000000;
12'd233 : tab2 = 23'b10110011011100100010010;
12'd234 : tab2 = 23'b10110011001010001110011;
12'd235 : tab2 = 23'b10110010110111111100000;
12'd236 : tab2 = 23'b10110010100101101010010;
12'd237 : tab2 = 23'b10110010010011011010000;
12'd238 : tab2 = 23'b10110010000001001011100;
12'd239 : tab2 = 23'b10110001101110111101101;
12'd240 : tab2 = 23'b10110001011100110001100;
12'd241 : tab2 = 23'b10110001001010100110010;
12'd242 : tab2 = 23'b10110000111000011100100;
12'd243 : tab2 = 23'b10110000100110010100000;
12'd244 : tab2 = 23'b10110000010100001100111;
12'd245 : tab2 = 23'b10110000000010000111000;
12'd246 : tab2 = 23'b10101111110000000010000;
12'd247 : tab2 = 23'b10101111011101111110100;
12'd248 : tab2 = 23'b10101111001011111100010;
12'd249 : tab2 = 23'b10101110111001111011010;
12'd250 : tab2 = 23'b10101110100111111100000;
12'd251 : tab2 = 23'b10101110010101111101010;
12'd252 : tab2 = 23'b10101110000100000000010;
12'd253 : tab2 = 23'b10101101110010000100000;
12'd254 : tab2 = 23'b10101101100000001001000;
12'd255 : tab2 = 23'b10101101001110001111111;
12'd256 : tab2 = 23'b10101100111100010111111;
12'd257 : tab2 = 23'b10101100101010100001000;
12'd258 : tab2 = 23'b10101100011000101011000;
12'd259 : tab2 = 23'b10101100000110110110100;
12'd260 : tab2 = 23'b10101011110101000010111;
12'd261 : tab2 = 23'b10101011100011010001000;
12'd262 : tab2 = 23'b10101011010001100000010;
12'd263 : tab2 = 23'b10101010111111110000110;
12'd264 : tab2 = 23'b10101010101110000010011;
12'd265 : tab2 = 23'b10101010011100010101011;
12'd266 : tab2 = 23'b10101010001010101001101;
12'd267 : tab2 = 23'b10101001111000111111000;
12'd268 : tab2 = 23'b10101001100111010101010;
12'd269 : tab2 = 23'b10101001010101101101010;
12'd270 : tab2 = 23'b10101001000100000110001;
12'd271 : tab2 = 23'b10101000110010100000001;
12'd272 : tab2 = 23'b10101000100000111100000;
12'd273 : tab2 = 23'b10101000001111011000010;
12'd274 : tab2 = 23'b10100111111101110110011;
12'd275 : tab2 = 23'b10100111101100010100111;
12'd276 : tab2 = 23'b10100111011010110101010;
12'd277 : tab2 = 23'b10100111001001010110110;
12'd278 : tab2 = 23'b10100110110111111001010;
12'd279 : tab2 = 23'b10100110100110011101010;
12'd280 : tab2 = 23'b10100110010101000010010;
12'd281 : tab2 = 23'b10100110000011101000011;
12'd282 : tab2 = 23'b10100101110010001111111;
12'd283 : tab2 = 23'b10100101100000111000100;
12'd284 : tab2 = 23'b10100101001111100010011;
12'd285 : tab2 = 23'b10100100111110001101011;
12'd286 : tab2 = 23'b10100100101100111001110;
12'd287 : tab2 = 23'b10100100011011100111000;
12'd288 : tab2 = 23'b10100100001010010101101;
12'd289 : tab2 = 23'b10100011111001000101001;
12'd290 : tab2 = 23'b10100011100111110110001;
12'd291 : tab2 = 23'b10100011010110101000010;
12'd292 : tab2 = 23'b10100011000101011011011;
12'd293 : tab2 = 23'b10100010110100010000000;
12'd294 : tab2 = 23'b10100010100011000101111;
12'd295 : tab2 = 23'b10100010010001111100011;
12'd296 : tab2 = 23'b10100010000000110100011;
12'd297 : tab2 = 23'b10100001101111101101101;
12'd298 : tab2 = 23'b10100001011110100111100;
12'd299 : tab2 = 23'b10100001001101100011010;
12'd300 : tab2 = 23'b10100000111100100000000;
12'd301 : tab2 = 23'b10100000101011011101101;
12'd302 : tab2 = 23'b10100000011010011100100;
12'd303 : tab2 = 23'b10100000001001011100111;
12'd304 : tab2 = 23'b10011111111000011110000;
12'd305 : tab2 = 23'b10011111100111100000101;
12'd306 : tab2 = 23'b10011111010110100100010;
12'd307 : tab2 = 23'b10011111000101101000111;
12'd308 : tab2 = 23'b10011110110100101110101;
12'd309 : tab2 = 23'b10011110100011110101111;
12'd310 : tab2 = 23'b10011110010010111101110;
12'd311 : tab2 = 23'b10011110000010000111010;
12'd312 : tab2 = 23'b10011101110001010001110;
12'd313 : tab2 = 23'b10011101100000011101011;
12'd314 : tab2 = 23'b10011101001111101010000;
12'd315 : tab2 = 23'b10011100111110110111101;
12'd316 : tab2 = 23'b10011100101110000110111;
12'd317 : tab2 = 23'b10011100011101010111010;
12'd318 : tab2 = 23'b10011100001100101000001;
12'd319 : tab2 = 23'b10011011111011111010101;
12'd320 : tab2 = 23'b10011011101011001110010;
12'd321 : tab2 = 23'b10011011011010100011001;
12'd322 : tab2 = 23'b10011011001001111001000;
12'd323 : tab2 = 23'b10011010111001001111011;
12'd324 : tab2 = 23'b10011010101000100111110;
12'd325 : tab2 = 23'b10011010011000000000100;
12'd326 : tab2 = 23'b10011010000111011010111;
12'd327 : tab2 = 23'b10011001110110110110100;
12'd328 : tab2 = 23'b10011001100110010010101;
12'd329 : tab2 = 23'b10011001010101110000110;
12'd330 : tab2 = 23'b10011001000101001111001;
12'd331 : tab2 = 23'b10011000110100101111001;
12'd332 : tab2 = 23'b10011000100100001111111;
12'd333 : tab2 = 23'b10011000010011110010001;
12'd334 : tab2 = 23'b10011000000011010101011;
12'd335 : tab2 = 23'b10010111110010111001101;
12'd336 : tab2 = 23'b10010111100010011110110;
12'd337 : tab2 = 23'b10010111010010000101101;
12'd338 : tab2 = 23'b10010111000001101100111;
12'd339 : tab2 = 23'b10010110110001010110000;
12'd340 : tab2 = 23'b10010110100000111111100;
12'd341 : tab2 = 23'b10010110010000101010011;
12'd342 : tab2 = 23'b10010110000000010110010;
12'd343 : tab2 = 23'b10010101110000000011000;
12'd344 : tab2 = 23'b10010101011111110001100;
12'd345 : tab2 = 23'b10010101001111100000011;
12'd346 : tab2 = 23'b10010100111111010000111;
12'd347 : tab2 = 23'b10010100101111000010101;
12'd348 : tab2 = 23'b10010100011110110100110;
12'd349 : tab2 = 23'b10010100001110101000010;
12'd350 : tab2 = 23'b10010011111110011100111;
12'd351 : tab2 = 23'b10010011101110010010110;
12'd352 : tab2 = 23'b10010011011110001001001;
12'd353 : tab2 = 23'b10010011001110000001011;
12'd354 : tab2 = 23'b10010010111101111010100;
12'd355 : tab2 = 23'b10010010101101110100110;
12'd356 : tab2 = 23'b10010010011101101111011;
12'd357 : tab2 = 23'b10010010001101101011100;
12'd358 : tab2 = 23'b10010001111101101000101;
12'd359 : tab2 = 23'b10010001101101100111001;
12'd360 : tab2 = 23'b10010001011101100110000;
12'd361 : tab2 = 23'b10010001001101100110101;
12'd362 : tab2 = 23'b10010000111101101000010;
12'd363 : tab2 = 23'b10010000101101101011001;
12'd364 : tab2 = 23'b10010000011101101110010;
12'd365 : tab2 = 23'b10010000001101110010100;
12'd366 : tab2 = 23'b10001111111101111000100;
12'd367 : tab2 = 23'b10001111101101111111100;
12'd368 : tab2 = 23'b10001111011110000111100;
12'd369 : tab2 = 23'b10001111001110010000011;
12'd370 : tab2 = 23'b10001110111110011010010;
12'd371 : tab2 = 23'b10001110101110100100110;
12'd372 : tab2 = 23'b10001110011110110001000;
12'd373 : tab2 = 23'b10001110001110111110011;
12'd374 : tab2 = 23'b10001101111111001100000;
12'd375 : tab2 = 23'b10001101101111011010111;
12'd376 : tab2 = 23'b10001101011111101011011;
12'd377 : tab2 = 23'b10001101001111111100101;
12'd378 : tab2 = 23'b10001101000000001111011;
12'd379 : tab2 = 23'b10001100110000100010001;
12'd380 : tab2 = 23'b10001100100000110110011;
12'd381 : tab2 = 23'b10001100010001001011100;
12'd382 : tab2 = 23'b10001100000001100010010;
12'd383 : tab2 = 23'b10001011110001111001111;
12'd384 : tab2 = 23'b10001011100010010010011;
12'd385 : tab2 = 23'b10001011010010101011100;
12'd386 : tab2 = 23'b10001011000011000101111;
12'd387 : tab2 = 23'b10001010110011100001100;
12'd388 : tab2 = 23'b10001010100011111110010;
12'd389 : tab2 = 23'b10001010010100011011101;
12'd390 : tab2 = 23'b10001010000100111010101;
12'd391 : tab2 = 23'b10001001110101011001111;
12'd392 : tab2 = 23'b10001001100101111010110;
12'd393 : tab2 = 23'b10001001010110011100010;
12'd394 : tab2 = 23'b10001001000110111110111;
12'd395 : tab2 = 23'b10001000110111100010100;
12'd396 : tab2 = 23'b10001000101000000111100;
12'd397 : tab2 = 23'b10001000011000101100111;
12'd398 : tab2 = 23'b10001000001001010011101;
12'd399 : tab2 = 23'b10000111111001111011011;
12'd400 : tab2 = 23'b10000111101010100100001;
12'd401 : tab2 = 23'b10000111011011001101101;
12'd402 : tab2 = 23'b10000111001011111000001;
12'd403 : tab2 = 23'b10000110111100100100000;
12'd404 : tab2 = 23'b10000110101101010000111;
12'd405 : tab2 = 23'b10000110011101111110100;
12'd406 : tab2 = 23'b10000110001110101101001;
12'd407 : tab2 = 23'b10000101111111011100110;
12'd408 : tab2 = 23'b10000101110000001101100;
12'd409 : tab2 = 23'b10000101100000111110111;
12'd410 : tab2 = 23'b10000101010001110001111;
12'd411 : tab2 = 23'b10000101000010100101010;
12'd412 : tab2 = 23'b10000100110011011001110;
12'd413 : tab2 = 23'b10000100100100001111111;
12'd414 : tab2 = 23'b10000100010101000110010;
12'd415 : tab2 = 23'b10000100000101111101111;
12'd416 : tab2 = 23'b10000011110110110110011;
12'd417 : tab2 = 23'b10000011100111110000010;
12'd418 : tab2 = 23'b10000011011000101010100;
12'd419 : tab2 = 23'b10000011001001100110000;
12'd420 : tab2 = 23'b10000010111010100010101;
12'd421 : tab2 = 23'b10000010101011100000001;
12'd422 : tab2 = 23'b10000010011100011110110;
12'd423 : tab2 = 23'b10000010001101011101110;
12'd424 : tab2 = 23'b10000001111110011110011;
12'd425 : tab2 = 23'b10000001101111100000000;
12'd426 : tab2 = 23'b10000001100000100010010;
12'd427 : tab2 = 23'b10000001010001100101001;
12'd428 : tab2 = 23'b10000001000010101001101;
12'd429 : tab2 = 23'b10000000110011101110110;
12'd430 : tab2 = 23'b10000000100100110100111;
12'd431 : tab2 = 23'b10000000010101111100001;
12'd432 : tab2 = 23'b10000000000111000100100;
12'd433 : tab2 = 23'b01111111111000001101010;
12'd434 : tab2 = 23'b01111111101001010111101;
12'd435 : tab2 = 23'b01111111011010100010011;
12'd436 : tab2 = 23'b01111111001011101110100;
12'd437 : tab2 = 23'b01111110111100111011001;
12'd438 : tab2 = 23'b01111110101110001001000;
12'd439 : tab2 = 23'b01111110011111011000000;
12'd440 : tab2 = 23'b01111110010000100111101;
12'd441 : tab2 = 23'b01111110000001111000010;
12'd442 : tab2 = 23'b01111101110011001001111;
12'd443 : tab2 = 23'b01111101100100011100101;
12'd444 : tab2 = 23'b01111101010101110000000;
12'd445 : tab2 = 23'b01111101000111000100011;
12'd446 : tab2 = 23'b01111100111000011001110;
12'd447 : tab2 = 23'b01111100101001110000010;
12'd448 : tab2 = 23'b01111100011011000111101;
12'd449 : tab2 = 23'b01111100001100011111110;
12'd450 : tab2 = 23'b01111011111101111000110;
12'd451 : tab2 = 23'b01111011101111010011001;
12'd452 : tab2 = 23'b01111011100000101110001;
12'd453 : tab2 = 23'b01111011010010001010001;
12'd454 : tab2 = 23'b01111011000011100110111;
12'd455 : tab2 = 23'b01111010110101000100110;
12'd456 : tab2 = 23'b01111010100110100011010;
12'd457 : tab2 = 23'b01111010011000000011001;
12'd458 : tab2 = 23'b01111010001001100100001;
12'd459 : tab2 = 23'b01111001111011000101100;
12'd460 : tab2 = 23'b01111001101100100111110;
12'd461 : tab2 = 23'b01111001011110001011010;
12'd462 : tab2 = 23'b01111001001111101111010;
12'd463 : tab2 = 23'b01111001000001010100100;
12'd464 : tab2 = 23'b01111000110010111010110;
12'd465 : tab2 = 23'b01111000100100100001111;
12'd466 : tab2 = 23'b01111000010110001001011;
12'd467 : tab2 = 23'b01111000000111110010111;
12'd468 : tab2 = 23'b01110111111001011100100;
12'd469 : tab2 = 23'b01110111101011000111100;
12'd470 : tab2 = 23'b01110111011100110010110;
12'd471 : tab2 = 23'b01110111001110011111011;
12'd472 : tab2 = 23'b01110111000000001100101;
12'd473 : tab2 = 23'b01110110110001111011010;
12'd474 : tab2 = 23'b01110110100011101010010;
12'd475 : tab2 = 23'b01110110010101011010010;
12'd476 : tab2 = 23'b01110110000111001011100;
12'd477 : tab2 = 23'b01110101111000111101111;
12'd478 : tab2 = 23'b01110101101010110000100;
12'd479 : tab2 = 23'b01110101011100100100001;
12'd480 : tab2 = 23'b01110101001110011001000;
12'd481 : tab2 = 23'b01110101000000001110001;
12'd482 : tab2 = 23'b01110100110010000101000;
12'd483 : tab2 = 23'b01110100100011111100001;
12'd484 : tab2 = 23'b01110100010101110100010;
12'd485 : tab2 = 23'b01110100000111101101010;
12'd486 : tab2 = 23'b01110011111001100111101;
12'd487 : tab2 = 23'b01110011101011100010011;
12'd488 : tab2 = 23'b01110011011101011110010;
12'd489 : tab2 = 23'b01110011001111011010111;
12'd490 : tab2 = 23'b01110011000001011000100;
12'd491 : tab2 = 23'b01110010110011010111000;
12'd492 : tab2 = 23'b01110010100101010110100;
12'd493 : tab2 = 23'b01110010010111010110101;
12'd494 : tab2 = 23'b01110010001001010111011;
12'd495 : tab2 = 23'b01110001111011011001010;
12'd496 : tab2 = 23'b01110001101101011100010;
12'd497 : tab2 = 23'b01110001011111100000001;
12'd498 : tab2 = 23'b01110001010001100100100;
12'd499 : tab2 = 23'b01110001000011101010100;
12'd500 : tab2 = 23'b01110000110101110000101;
12'd501 : tab2 = 23'b01110000100111110111100;
12'd502 : tab2 = 23'b01110000011001111111111;
12'd503 : tab2 = 23'b01110000001100001000110;
12'd504 : tab2 = 23'b01101111111110010010100;
12'd505 : tab2 = 23'b01101111110000011101100;
12'd506 : tab2 = 23'b01101111100010101000110;
12'd507 : tab2 = 23'b01101111010100110101101;
12'd508 : tab2 = 23'b01101111000111000010111;
12'd509 : tab2 = 23'b01101110111001010000110;
12'd510 : tab2 = 23'b01101110101011011111111;
12'd511 : tab2 = 23'b01101110011101101111111;
12'd512 : tab2 = 23'b01101110010000000000101;
12'd513 : tab2 = 23'b01101110000010010010010;
12'd514 : tab2 = 23'b01101101110100100100010;
12'd515 : tab2 = 23'b01101101100110110111110;
12'd516 : tab2 = 23'b01101101011001001100010;
12'd517 : tab2 = 23'b01101101001011100001000;
12'd518 : tab2 = 23'b01101100111101110110111;
12'd519 : tab2 = 23'b01101100110000001101110;
12'd520 : tab2 = 23'b01101100100010100101001;
12'd521 : tab2 = 23'b01101100010100111110000;
12'd522 : tab2 = 23'b01101100000111010111001;
12'd523 : tab2 = 23'b01101011111001110001000;
12'd524 : tab2 = 23'b01101011101100001011110;
12'd525 : tab2 = 23'b01101011011110100111110;
12'd526 : tab2 = 23'b01101011010001000100011;
12'd527 : tab2 = 23'b01101011000011100010000;
12'd528 : tab2 = 23'b01101010110110000000010;
12'd529 : tab2 = 23'b01101010101000011111011;
12'd530 : tab2 = 23'b01101010011010111111011;
12'd531 : tab2 = 23'b01101010001101100000100;
12'd532 : tab2 = 23'b01101010000000000010011;
12'd533 : tab2 = 23'b01101001110010100100011;
12'd534 : tab2 = 23'b01101001100101000111111;
12'd535 : tab2 = 23'b01101001010111101100000;
12'd536 : tab2 = 23'b01101001001010010001000;
12'd537 : tab2 = 23'b01101000111100110110110;
12'd538 : tab2 = 23'b01101000101111011101011;
12'd539 : tab2 = 23'b01101000100010000101001;
12'd540 : tab2 = 23'b01101000010100101101010;
12'd541 : tab2 = 23'b01101000000111010110011;
12'd542 : tab2 = 23'b01100111111010000000011;
12'd543 : tab2 = 23'b01100111101100101011010;
12'd544 : tab2 = 23'b01100111011111010110111;
12'd545 : tab2 = 23'b01100111010010000011011;
12'd546 : tab2 = 23'b01100111000100110000110;
12'd547 : tab2 = 23'b01100110110111011110011;
12'd548 : tab2 = 23'b01100110101010001101110;
12'd549 : tab2 = 23'b01100110011100111101010;
12'd550 : tab2 = 23'b01100110001111101110000;
12'd551 : tab2 = 23'b01100110000010011111001;
12'd552 : tab2 = 23'b01100101110101010001110;
12'd553 : tab2 = 23'b01100101101000000100110;
12'd554 : tab2 = 23'b01100101011010111000010;
12'd555 : tab2 = 23'b01100101001101101100110;
12'd556 : tab2 = 23'b01100101000000100010001;
12'd557 : tab2 = 23'b01100100110011011000011;
12'd558 : tab2 = 23'b01100100100110001111011;
12'd559 : tab2 = 23'b01100100011001000111001;
12'd560 : tab2 = 23'b01100100001011111111111;
12'd561 : tab2 = 23'b01100011111110111001101;
12'd562 : tab2 = 23'b01100011110001110011111;
12'd563 : tab2 = 23'b01100011100100101110111;
12'd564 : tab2 = 23'b01100011010111101010110;
12'd565 : tab2 = 23'b01100011001010100111100;
12'd566 : tab2 = 23'b01100010111101100101000;
12'd567 : tab2 = 23'b01100010110000100010111;
12'd568 : tab2 = 23'b01100010100011100010011;
12'd569 : tab2 = 23'b01100010010110100001110;
12'd570 : tab2 = 23'b01100010001001100010110;
12'd571 : tab2 = 23'b01100001111100100011110;
12'd572 : tab2 = 23'b01100001101111100110001;
12'd573 : tab2 = 23'b01100001100010101001001;
12'd574 : tab2 = 23'b01100001010101101101001;
12'd575 : tab2 = 23'b01100001001000110001101;
12'd576 : tab2 = 23'b01100000111011110110111;
12'd577 : tab2 = 23'b01100000101110111101000;
12'd578 : tab2 = 23'b01100000100010000100010;
12'd579 : tab2 = 23'b01100000010101001011110;
12'd580 : tab2 = 23'b01100000001000010100010;
12'd581 : tab2 = 23'b01011111111011011101101;
12'd582 : tab2 = 23'b01011111101110100111101;
12'd583 : tab2 = 23'b01011111100001110010100;
12'd584 : tab2 = 23'b01011111010100111110010;
12'd585 : tab2 = 23'b01011111001000001010111;
12'd586 : tab2 = 23'b01011110111011010111111;
12'd587 : tab2 = 23'b01011110101110100101110;
12'd588 : tab2 = 23'b01011110100001110100111;
12'd589 : tab2 = 23'b01011110010101000100010;
12'd590 : tab2 = 23'b01011110001000010100100;
12'd591 : tab2 = 23'b01011101111011100101010;
12'd592 : tab2 = 23'b01011101101110110111010;
12'd593 : tab2 = 23'b01011101100010001010000;
12'd594 : tab2 = 23'b01011101010101011101001;
12'd595 : tab2 = 23'b01011101001000110001011;
12'd596 : tab2 = 23'b01011100111100000110010;
12'd597 : tab2 = 23'b01011100101111011100010;
12'd598 : tab2 = 23'b01011100100010110010110;
12'd599 : tab2 = 23'b01011100010110001001100;
12'd600 : tab2 = 23'b01011100001001100001100;
12'd601 : tab2 = 23'b01011011111100111010011;
12'd602 : tab2 = 23'b01011011110000010100001;
12'd603 : tab2 = 23'b01011011100011101110001;
12'd604 : tab2 = 23'b01011011010111001001000;
12'd605 : tab2 = 23'b01011011001010100100111;
12'd606 : tab2 = 23'b01011010111110000001101;
12'd607 : tab2 = 23'b01011010110001011110111;
12'd608 : tab2 = 23'b01011010100100111101000;
12'd609 : tab2 = 23'b01011010011000011011110;
12'd610 : tab2 = 23'b01011010001011111011100;
12'd611 : tab2 = 23'b01011001111111011011110;
12'd612 : tab2 = 23'b01011001110010111100110;
12'd613 : tab2 = 23'b01011001100110011110100;
12'd614 : tab2 = 23'b01011001011010000001000;
12'd615 : tab2 = 23'b01011001001101100100100;
12'd616 : tab2 = 23'b01011001000001001000100;
12'd617 : tab2 = 23'b01011000110100101101100;
12'd618 : tab2 = 23'b01011000101000010010111;
12'd619 : tab2 = 23'b01011000011011111000101;
12'd620 : tab2 = 23'b01011000001111100000000;
12'd621 : tab2 = 23'b01011000000011001000000;
12'd622 : tab2 = 23'b01010111110110110000100;
12'd623 : tab2 = 23'b01010111101010011001110;
12'd624 : tab2 = 23'b01010111011110000011101;
12'd625 : tab2 = 23'b01010111010001101110011;
12'd626 : tab2 = 23'b01010111000101011001110;
12'd627 : tab2 = 23'b01010110111001000101111;
12'd628 : tab2 = 23'b01010110101100110011000;
12'd629 : tab2 = 23'b01010110100000100000111;
12'd630 : tab2 = 23'b01010110010100001111001;
12'd631 : tab2 = 23'b01010110000111111110001;
12'd632 : tab2 = 23'b01010101111011101110001;
12'd633 : tab2 = 23'b01010101101111011110101;
12'd634 : tab2 = 23'b01010101100011010000001;
12'd635 : tab2 = 23'b01010101010111000010101;
12'd636 : tab2 = 23'b01010101001010110100111;
12'd637 : tab2 = 23'b01010100111110101000100;
12'd638 : tab2 = 23'b01010100110010011100100;
12'd639 : tab2 = 23'b01010100100110010010000;
12'd640 : tab2 = 23'b01010100011010000111100;
12'd641 : tab2 = 23'b01010100001101111110000;
12'd642 : tab2 = 23'b01010100000001110101001;
12'd643 : tab2 = 23'b01010011110101101101001;
12'd644 : tab2 = 23'b01010011101001100101100;
12'd645 : tab2 = 23'b01010011011101011110111;
12'd646 : tab2 = 23'b01010011010001011000101;
12'd647 : tab2 = 23'b01010011000101010011111;
12'd648 : tab2 = 23'b01010010111001001111010;
12'd649 : tab2 = 23'b01010010101101001011100;
12'd650 : tab2 = 23'b01010010100001001000001;
12'd651 : tab2 = 23'b01010010010101000101111;
12'd652 : tab2 = 23'b01010010001001000011111;
12'd653 : tab2 = 23'b01010001111101000010111;
12'd654 : tab2 = 23'b01010001110001000011000;
12'd655 : tab2 = 23'b01010001100101000011101;
12'd656 : tab2 = 23'b01010001011001000100011;
12'd657 : tab2 = 23'b01010001001101000110011;
12'd658 : tab2 = 23'b01010001000001001000111;
12'd659 : tab2 = 23'b01010000110101001100011;
12'd660 : tab2 = 23'b01010000101001010000011;
12'd661 : tab2 = 23'b01010000011101010101001;
12'd662 : tab2 = 23'b01010000010001011010010;
12'd663 : tab2 = 23'b01010000000101100000110;
12'd664 : tab2 = 23'b01001111111001100111010;
12'd665 : tab2 = 23'b01001111101101101111001;
12'd666 : tab2 = 23'b01001111100001110111001;
12'd667 : tab2 = 23'b01001111010101111111111;
12'd668 : tab2 = 23'b01001111001010001001100;
12'd669 : tab2 = 23'b01001110111110010100000;
12'd670 : tab2 = 23'b01001110110010011111010;
12'd671 : tab2 = 23'b01001110100110101010101;
12'd672 : tab2 = 23'b01001110011010110111000;
12'd673 : tab2 = 23'b01001110001111000100000;
12'd674 : tab2 = 23'b01001110000011010010001;
12'd675 : tab2 = 23'b01001101110111100000100;
12'd676 : tab2 = 23'b01001101101011101111110;
12'd677 : tab2 = 23'b01001101011111111111110;
12'd678 : tab2 = 23'b01001101010100010000001;
12'd679 : tab2 = 23'b01001101001000100001010;
12'd680 : tab2 = 23'b01001100111100110011010;
12'd681 : tab2 = 23'b01001100110001000101100;
12'd682 : tab2 = 23'b01001100100101011001000;
12'd683 : tab2 = 23'b01001100011001101101010;
12'd684 : tab2 = 23'b01001100001110000001110;
12'd685 : tab2 = 23'b01001100000010010111001;
12'd686 : tab2 = 23'b01001011110110101101010;
12'd687 : tab2 = 23'b01001011101011000011110;
12'd688 : tab2 = 23'b01001011011111011011011;
12'd689 : tab2 = 23'b01001011010011110011001;
12'd690 : tab2 = 23'b01001011001000001011111;
12'd691 : tab2 = 23'b01001010111100100101011;
12'd692 : tab2 = 23'b01001010110000111111100;
12'd693 : tab2 = 23'b01001010100101011010011;
12'd694 : tab2 = 23'b01001010011001110101110;
12'd695 : tab2 = 23'b01001010001110010010000;
12'd696 : tab2 = 23'b01001010000010101110101;
12'd697 : tab2 = 23'b01001001110111001100011;
12'd698 : tab2 = 23'b01001001101011101010001;
12'd699 : tab2 = 23'b01001001100000001001010;
12'd700 : tab2 = 23'b01001001010100101000100;
12'd701 : tab2 = 23'b01001001001001001001000;
12'd702 : tab2 = 23'b01001000111101101001101;
12'd703 : tab2 = 23'b01001000110010001011011;
12'd704 : tab2 = 23'b01001000100110101101011;
12'd705 : tab2 = 23'b01001000011011010000011;
12'd706 : tab2 = 23'b01001000001111110011100;
12'd707 : tab2 = 23'b01001000000100010111110;
12'd708 : tab2 = 23'b01000111111000111100110;
12'd709 : tab2 = 23'b01000111101101100010011;
12'd710 : tab2 = 23'b01000111100010001000010;
12'd711 : tab2 = 23'b01000111010110101111001;
12'd712 : tab2 = 23'b01000111001011010110110;
12'd713 : tab2 = 23'b01000110111111111110110;
12'd714 : tab2 = 23'b01000110110100100111110;
12'd715 : tab2 = 23'b01000110101001010001011;
12'd716 : tab2 = 23'b01000110011101111011000;
12'd717 : tab2 = 23'b01000110010010100110001;
12'd718 : tab2 = 23'b01000110000111010001011;
12'd719 : tab2 = 23'b01000101111011111101101;
12'd720 : tab2 = 23'b01000101110000101001111;
12'd721 : tab2 = 23'b01000101100101010111011;
12'd722 : tab2 = 23'b01000101011010000101011;
12'd723 : tab2 = 23'b01000101001110110100000;
12'd724 : tab2 = 23'b01000101000011100011101;
12'd725 : tab2 = 23'b01000100111000010011100;
12'd726 : tab2 = 23'b01000100101101000100000;
12'd727 : tab2 = 23'b01000100100001110101100;
12'd728 : tab2 = 23'b01000100010110100111101;
12'd729 : tab2 = 23'b01000100001011011010010;
12'd730 : tab2 = 23'b01000100000000001101001;
12'd731 : tab2 = 23'b01000011110101000001000;
12'd732 : tab2 = 23'b01000011101001110101111;
12'd733 : tab2 = 23'b01000011011110101010101;
12'd734 : tab2 = 23'b01000011010011100000011;
12'd735 : tab2 = 23'b01000011001000010111000;
12'd736 : tab2 = 23'b01000010111101001110010;
12'd737 : tab2 = 23'b01000010110010000101101;
12'd738 : tab2 = 23'b01000010100110111101111;
12'd739 : tab2 = 23'b01000010011011110110111;
12'd740 : tab2 = 23'b01000010010000110000110;
12'd741 : tab2 = 23'b01000010000101101010111;
12'd742 : tab2 = 23'b01000001111010100101110;
12'd743 : tab2 = 23'b01000001101111100001100;
12'd744 : tab2 = 23'b01000001100100011101100;
12'd745 : tab2 = 23'b01000001011001011010100;
12'd746 : tab2 = 23'b01000001001110010111110;
12'd747 : tab2 = 23'b01000001000011010110001;
12'd748 : tab2 = 23'b01000000111000010100100;
12'd749 : tab2 = 23'b01000000101101010100010;
12'd750 : tab2 = 23'b01000000100010010011111;
12'd751 : tab2 = 23'b01000000010111010100011;
12'd752 : tab2 = 23'b01000000001100010101110;
12'd753 : tab2 = 23'b01000000000001010111110;
12'd754 : tab2 = 23'b00111111110110011010000;
12'd755 : tab2 = 23'b00111111101011011101000;
12'd756 : tab2 = 23'b00111111100000100000111;
12'd757 : tab2 = 23'b00111111010101100101010;
12'd758 : tab2 = 23'b00111111001010101010011;
12'd759 : tab2 = 23'b00111110111111101111110;
12'd760 : tab2 = 23'b00111110110100110110001;
12'd761 : tab2 = 23'b00111110101001111100111;
12'd762 : tab2 = 23'b00111110011111000100010;
12'd763 : tab2 = 23'b00111110010100001100011;
12'd764 : tab2 = 23'b00111110001001010101000;
12'd765 : tab2 = 23'b00111101111110011110011;
12'd766 : tab2 = 23'b00111101110011101000001;
12'd767 : tab2 = 23'b00111101101000110010111;
12'd768 : tab2 = 23'b00111101011101111101111;
12'd769 : tab2 = 23'b00111101010011001001101;
12'd770 : tab2 = 23'b00111101001000010110010;
12'd771 : tab2 = 23'b00111100111101100011010;
12'd772 : tab2 = 23'b00111100110010110001000;
12'd773 : tab2 = 23'b00111100100111111110111;
12'd774 : tab2 = 23'b00111100011101001101110;
12'd775 : tab2 = 23'b00111100010010011101001;
12'd776 : tab2 = 23'b00111100000111101101011;
12'd777 : tab2 = 23'b00111011111100111110001;
12'd778 : tab2 = 23'b00111011110010001111001;
12'd779 : tab2 = 23'b00111011100111100000111;
12'd780 : tab2 = 23'b00111011011100110011100;
12'd781 : tab2 = 23'b00111011010010000110100;
12'd782 : tab2 = 23'b00111011000111011010011;
12'd783 : tab2 = 23'b00111010111100101110110;
12'd784 : tab2 = 23'b00111010110010000011011;
12'd785 : tab2 = 23'b00111010100111011001010;
12'd786 : tab2 = 23'b00111010011100101111010;
12'd787 : tab2 = 23'b00111010010010000101111;
12'd788 : tab2 = 23'b00111010000111011101001;
12'd789 : tab2 = 23'b00111001111100110101001;
12'd790 : tab2 = 23'b00111001110010001101100;
12'd791 : tab2 = 23'b00111001100111100110110;
12'd792 : tab2 = 23'b00111001011101000000011;
12'd793 : tab2 = 23'b00111001010010011010101;
12'd794 : tab2 = 23'b00111001000111110101011;
12'd795 : tab2 = 23'b00111000111101010001000;
12'd796 : tab2 = 23'b00111000110010101101011;
12'd797 : tab2 = 23'b00111000101000001001101;
12'd798 : tab2 = 23'b00111000011101100111010;
12'd799 : tab2 = 23'b00111000010011000101000;
12'd800 : tab2 = 23'b00111000001000100011101;
12'd801 : tab2 = 23'b00110111111110000010100;
12'd802 : tab2 = 23'b00110111110011100001111;
12'd803 : tab2 = 23'b00110111101001000010010;
12'd804 : tab2 = 23'b00110111011110100011010;
12'd805 : tab2 = 23'b00110111010100000100110;
12'd806 : tab2 = 23'b00110111001001100110101;
12'd807 : tab2 = 23'b00110110111111001000111;
12'd808 : tab2 = 23'b00110110110100101100011;
12'd809 : tab2 = 23'b00110110101010010000000;
12'd810 : tab2 = 23'b00110110011111110100101;
12'd811 : tab2 = 23'b00110110010101011001010;
12'd812 : tab2 = 23'b00110110001010111110110;
12'd813 : tab2 = 23'b00110110000000100100100;
12'd814 : tab2 = 23'b00110101110110001011101;
12'd815 : tab2 = 23'b00110101101011110010110;
12'd816 : tab2 = 23'b00110101100001011010101;
12'd817 : tab2 = 23'b00110101010111000011001;
12'd818 : tab2 = 23'b00110101001100101100000;
12'd819 : tab2 = 23'b00110101000010010101100;
12'd820 : tab2 = 23'b00110100110111111111101;
12'd821 : tab2 = 23'b00110100101101101010011;
12'd822 : tab2 = 23'b00110100100011010101101;
12'd823 : tab2 = 23'b00110100011001000001110;
12'd824 : tab2 = 23'b00110100001110101110000;
12'd825 : tab2 = 23'b00110100000100011011000;
12'd826 : tab2 = 23'b00110011111010001000101;
12'd827 : tab2 = 23'b00110011101111110110110;
12'd828 : tab2 = 23'b00110011100101100101100;
12'd829 : tab2 = 23'b00110011011011010100111;
12'd830 : tab2 = 23'b00110011010001000100011;
12'd831 : tab2 = 23'b00110011000110110101010;
12'd832 : tab2 = 23'b00110010111100100110011;
12'd833 : tab2 = 23'b00110010110010010111111;
12'd834 : tab2 = 23'b00110010101000001001101;
12'd835 : tab2 = 23'b00110010011101111100100;
12'd836 : tab2 = 23'b00110010010011110000001;
12'd837 : tab2 = 23'b00110010001001100011100;
12'd838 : tab2 = 23'b00110001111111011000001;
12'd839 : tab2 = 23'b00110001110101001101001;
12'd840 : tab2 = 23'b00110001101011000010101;
12'd841 : tab2 = 23'b00110001100000111000110;
12'd842 : tab2 = 23'b00110001010110101111010;
12'd843 : tab2 = 23'b00110001001100100110010;
12'd844 : tab2 = 23'b00110001000010011110011;
12'd845 : tab2 = 23'b00110000111000010110101;
12'd846 : tab2 = 23'b00110000101110001111101;
12'd847 : tab2 = 23'b00110000100100001001000;
12'd848 : tab2 = 23'b00110000011010000011000;
12'd849 : tab2 = 23'b00110000001111111101101;
12'd850 : tab2 = 23'b00110000000101111001001;
12'd851 : tab2 = 23'b00101111111011110100010;
12'd852 : tab2 = 23'b00101111110001110000110;
12'd853 : tab2 = 23'b00101111100111101101101;
12'd854 : tab2 = 23'b00101111011101101010111;
12'd855 : tab2 = 23'b00101111010011101000110;
12'd856 : tab2 = 23'b00101111001001100111011;
12'd857 : tab2 = 23'b00101110111111100110000;
12'd858 : tab2 = 23'b00101110110101100110000;
12'd859 : tab2 = 23'b00101110101011100101111;
12'd860 : tab2 = 23'b00101110100001100110100;
12'd861 : tab2 = 23'b00101110010111100111110;
12'd862 : tab2 = 23'b00101110001101101001101;
12'd863 : tab2 = 23'b00101110000011101100000;
12'd864 : tab2 = 23'b00101101111001101110110;
12'd865 : tab2 = 23'b00101101101111110010001;
12'd866 : tab2 = 23'b00101101100101110110001;
12'd867 : tab2 = 23'b00101101011011111010101;
12'd868 : tab2 = 23'b00101101010001111111101;
12'd869 : tab2 = 23'b00101101001000000101011;
12'd870 : tab2 = 23'b00101100111110001011110;
12'd871 : tab2 = 23'b00101100110100010001111;
12'd872 : tab2 = 23'b00101100101010011001011;
12'd873 : tab2 = 23'b00101100100000100001010;
12'd874 : tab2 = 23'b00101100010110101001001;
12'd875 : tab2 = 23'b00101100001100110010010;
12'd876 : tab2 = 23'b00101100000010111011011;
12'd877 : tab2 = 23'b00101011111001000101100;
12'd878 : tab2 = 23'b00101011101111001111110;
12'd879 : tab2 = 23'b00101011100101011010101;
12'd880 : tab2 = 23'b00101011011011100110011;
12'd881 : tab2 = 23'b00101011010001110010001;
12'd882 : tab2 = 23'b00101011000111111110111;
12'd883 : tab2 = 23'b00101010111110001100001;
12'd884 : tab2 = 23'b00101010110100011001111;
12'd885 : tab2 = 23'b00101010101010101000011;
12'd886 : tab2 = 23'b00101010100000110110110;
12'd887 : tab2 = 23'b00101010010111000101110;
12'd888 : tab2 = 23'b00101010001101010101110;
12'd889 : tab2 = 23'b00101010000011100101110;
12'd890 : tab2 = 23'b00101001111001110110111;
12'd891 : tab2 = 23'b00101001110000001000011;
12'd892 : tab2 = 23'b00101001100110011010100;
12'd893 : tab2 = 23'b00101001011100101100110;
12'd894 : tab2 = 23'b00101001010010111111101;
12'd895 : tab2 = 23'b00101001001001010011000;
12'd896 : tab2 = 23'b00101000111111100111010;
12'd897 : tab2 = 23'b00101000110101111011101;
12'd898 : tab2 = 23'b00101000101100010000110;
12'd899 : tab2 = 23'b00101000100010100110011;
12'd900 : tab2 = 23'b00101000011000111100110;
12'd901 : tab2 = 23'b00101000001111010011010;
12'd902 : tab2 = 23'b00101000000101101010011;
12'd903 : tab2 = 23'b00100111111100000010010;
12'd904 : tab2 = 23'b00100111110010011010001;
12'd905 : tab2 = 23'b00100111101000110011011;
12'd906 : tab2 = 23'b00100111011111001100010;
12'd907 : tab2 = 23'b00100111010101100110010;
12'd908 : tab2 = 23'b00100111001100000000000;
12'd909 : tab2 = 23'b00100111000010011011001;
12'd910 : tab2 = 23'b00100110111000110110011;
12'd911 : tab2 = 23'b00100110101111010010011;
12'd912 : tab2 = 23'b00100110100101101110110;
12'd913 : tab2 = 23'b00100110011100001011110;
12'd914 : tab2 = 23'b00100110010010101001001;
12'd915 : tab2 = 23'b00100110001001000111000;
12'd916 : tab2 = 23'b00100101111111100101010;
12'd917 : tab2 = 23'b00100101110110000100011;
12'd918 : tab2 = 23'b00100101101100100011111;
12'd919 : tab2 = 23'b00100101100011000011101;
12'd920 : tab2 = 23'b00100101011001100100010;
12'd921 : tab2 = 23'b00100101010000000101001;
12'd922 : tab2 = 23'b00100101000110100110110;
12'd923 : tab2 = 23'b00100100111101001001001;
12'd924 : tab2 = 23'b00100100110011101011011;
12'd925 : tab2 = 23'b00100100101010001110011;
12'd926 : tab2 = 23'b00100100100000110010001;
12'd927 : tab2 = 23'b00100100010111010110000;
12'd928 : tab2 = 23'b00100100001101111010101;
12'd929 : tab2 = 23'b00100100000100011111100;
12'd930 : tab2 = 23'b00100011111011000101000;
12'd931 : tab2 = 23'b00100011110001101011011;
12'd932 : tab2 = 23'b00100011101000010001111;
12'd933 : tab2 = 23'b00100011011110111001000;
12'd934 : tab2 = 23'b00100011010101100000100;
12'd935 : tab2 = 23'b00100011001100001000101;
12'd936 : tab2 = 23'b00100011000010110001100;
12'd937 : tab2 = 23'b00100010111001011010100;
12'd938 : tab2 = 23'b00100010110000000100000;
12'd939 : tab2 = 23'b00100010100110101110000;
12'd940 : tab2 = 23'b00100010011101011000011;
12'd941 : tab2 = 23'b00100010010100000011110;
12'd942 : tab2 = 23'b00100010001010101111010;
12'd943 : tab2 = 23'b00100010000001011011010;
12'd944 : tab2 = 23'b00100001111000001000000;
12'd945 : tab2 = 23'b00100001101110110101001;
12'd946 : tab2 = 23'b00100001100101100010101;
12'd947 : tab2 = 23'b00100001011100010000111;
12'd948 : tab2 = 23'b00100001010010111111011;
12'd949 : tab2 = 23'b00100001001001101110011;
12'd950 : tab2 = 23'b00100001000000011101111;
12'd951 : tab2 = 23'b00100000110111001110011;
12'd952 : tab2 = 23'b00100000101101111110110;
12'd953 : tab2 = 23'b00100000100100101111110;
12'd954 : tab2 = 23'b00100000011011100001010;
12'd955 : tab2 = 23'b00100000010010010011000;
12'd956 : tab2 = 23'b00100000001001000101110;
12'd957 : tab2 = 23'b00011111111111111000101;
12'd958 : tab2 = 23'b00011111110110101100010;
12'd959 : tab2 = 23'b00011111101101100000011;
12'd960 : tab2 = 23'b00011111100100010100101;
12'd961 : tab2 = 23'b00011111011011001001110;
12'd962 : tab2 = 23'b00011111010001111111010;
12'd963 : tab2 = 23'b00011111001000110101001;
12'd964 : tab2 = 23'b00011110111111101011011;
12'd965 : tab2 = 23'b00011110110110100010101;
12'd966 : tab2 = 23'b00011110101101011001111;
12'd967 : tab2 = 23'b00011110100100010001110;
12'd968 : tab2 = 23'b00011110011011001010001;
12'd969 : tab2 = 23'b00011110010010000010111;
12'd970 : tab2 = 23'b00011110001000111100100;
12'd971 : tab2 = 23'b00011101111111110110011;
12'd972 : tab2 = 23'b00011101110110110000010;
12'd973 : tab2 = 23'b00011101101101101011100;
12'd974 : tab2 = 23'b00011101100100100110100;
12'd975 : tab2 = 23'b00011101011011100010010;
12'd976 : tab2 = 23'b00011101010010011110011;
12'd977 : tab2 = 23'b00011101001001011011011;
12'd978 : tab2 = 23'b00011101000000011000011;
12'd979 : tab2 = 23'b00011100110111010101111;
12'd980 : tab2 = 23'b00011100101110010100001;
12'd981 : tab2 = 23'b00011100100101010010110;
12'd982 : tab2 = 23'b00011100011100010001111;
12'd983 : tab2 = 23'b00011100010011010001010;
12'd984 : tab2 = 23'b00011100001010010001001;
12'd985 : tab2 = 23'b00011100000001010001111;
12'd986 : tab2 = 23'b00011011111000010010110;
12'd987 : tab2 = 23'b00011011101111010100011;
12'd988 : tab2 = 23'b00011011100110010110001;
12'd989 : tab2 = 23'b00011011011101011000111;
12'd990 : tab2 = 23'b00011011010100011011110;
12'd991 : tab2 = 23'b00011011001011011110111;
12'd992 : tab2 = 23'b00011011000010100010101;
12'd993 : tab2 = 23'b00011010111001100111010;
12'd994 : tab2 = 23'b00011010110000101011111;
12'd995 : tab2 = 23'b00011010100111110001000;
12'd996 : tab2 = 23'b00011010011110110110110;
12'd997 : tab2 = 23'b00011010010101111101000;
12'd998 : tab2 = 23'b00011010001101000011101;
12'd999 : tab2 = 23'b00011010000100001010110;
12'd1000 : tab2 = 23'b00011001111011010010010;
12'd1001 : tab2 = 23'b00011001110010011010010;
12'd1002 : tab2 = 23'b00011001101001100011000;
12'd1003 : tab2 = 23'b00011001100000101011101;
12'd1004 : tab2 = 23'b00011001010111110101010;
12'd1005 : tab2 = 23'b00011001001110111110111;
12'd1006 : tab2 = 23'b00011001000110001001001;
12'd1007 : tab2 = 23'b00011000111101010100010;
12'd1008 : tab2 = 23'b00011000110100011111010;
12'd1009 : tab2 = 23'b00011000101011101011010;
12'd1010 : tab2 = 23'b00011000100010110111100;
12'd1011 : tab2 = 23'b00011000011010000100011;
12'd1012 : tab2 = 23'b00011000010001010001001;
12'd1013 : tab2 = 23'b00011000001000011110101;
12'd1014 : tab2 = 23'b00010111111111101100111;
12'd1015 : tab2 = 23'b00010111110110111011011;
12'd1016 : tab2 = 23'b00010111101110001010100;
12'd1017 : tab2 = 23'b00010111100101011001101;
12'd1018 : tab2 = 23'b00010111011100101001010;
12'd1019 : tab2 = 23'b00010111010011111001111;
12'd1020 : tab2 = 23'b00010111001011001010110;
12'd1021 : tab2 = 23'b00010111000010011100001;
12'd1022 : tab2 = 23'b00010110111001101101101;
12'd1023 : tab2 = 23'b00010110110000111111111;
12'd1024 : tab2 = 23'b00010110101000010010011;
12'd1025 : tab2 = 23'b00010110011111100101010;
12'd1026 : tab2 = 23'b00010110010110111001010;
12'd1027 : tab2 = 23'b00010110001110001101000;
12'd1028 : tab2 = 23'b00010110000101100001100;
12'd1029 : tab2 = 23'b00010101111100110110011;
12'd1030 : tab2 = 23'b00010101110100001011100;
12'd1031 : tab2 = 23'b00010101101011100001001;
12'd1032 : tab2 = 23'b00010101100010110111101;
12'd1033 : tab2 = 23'b00010101011010001110010;
12'd1034 : tab2 = 23'b00010101010001100101010;
12'd1035 : tab2 = 23'b00010101001000111101000;
12'd1036 : tab2 = 23'b00010101000000010100111;
12'd1037 : tab2 = 23'b00010100110111101101100;
12'd1038 : tab2 = 23'b00010100101111000110010;
12'd1039 : tab2 = 23'b00010100100110011111101;
12'd1040 : tab2 = 23'b00010100011101111001101;
12'd1041 : tab2 = 23'b00010100010101010011101;
12'd1042 : tab2 = 23'b00010100001100101110011;
12'd1043 : tab2 = 23'b00010100000100001001100;
12'd1044 : tab2 = 23'b00010011111011100101010;
12'd1045 : tab2 = 23'b00010011110011000001000;
12'd1046 : tab2 = 23'b00010011101010011101100;
12'd1047 : tab2 = 23'b00010011100001111010101;
12'd1048 : tab2 = 23'b00010011011001010111111;
12'd1049 : tab2 = 23'b00010011010000110101100;
12'd1050 : tab2 = 23'b00010011001000010011111;
12'd1051 : tab2 = 23'b00010010111111110010110;
12'd1052 : tab2 = 23'b00010010110111010001011;
12'd1053 : tab2 = 23'b00010010101110110001000;
12'd1054 : tab2 = 23'b00010010100110010001001;
12'd1055 : tab2 = 23'b00010010011101110001101;
12'd1056 : tab2 = 23'b00010010010101010010010;
12'd1057 : tab2 = 23'b00010010001100110011101;
12'd1058 : tab2 = 23'b00010010000100010101101;
12'd1059 : tab2 = 23'b00010001111011110111100;
12'd1060 : tab2 = 23'b00010001110011011010001;
12'd1061 : tab2 = 23'b00010001101010111101001;
12'd1062 : tab2 = 23'b00010001100010100000110;
12'd1063 : tab2 = 23'b00010001011010000100101;
12'd1064 : tab2 = 23'b00010001010001101000101;
12'd1065 : tab2 = 23'b00010001001001001101101;
12'd1066 : tab2 = 23'b00010001000000110010110;
12'd1067 : tab2 = 23'b00010000111000011000100;
12'd1068 : tab2 = 23'b00010000101111111110110;
12'd1069 : tab2 = 23'b00010000100111100101011;
12'd1070 : tab2 = 23'b00010000011111001100001;
12'd1071 : tab2 = 23'b00010000010110110011100;
12'd1072 : tab2 = 23'b00010000001110011011100;
12'd1073 : tab2 = 23'b00010000000110000011101;
12'd1074 : tab2 = 23'b00001111111101101100010;
12'd1075 : tab2 = 23'b00001111110101010101001;
12'd1076 : tab2 = 23'b00001111101100111110101;
12'd1077 : tab2 = 23'b00001111100100101000111;
12'd1078 : tab2 = 23'b00001111011100010011010;
12'd1079 : tab2 = 23'b00001111010011111101111;
12'd1080 : tab2 = 23'b00001111001011101001000;
12'd1081 : tab2 = 23'b00001111000011010100111;
12'd1082 : tab2 = 23'b00001110111011000000101;
12'd1083 : tab2 = 23'b00001110110010101101100;
12'd1084 : tab2 = 23'b00001110101010011010000;
12'd1085 : tab2 = 23'b00001110100010000111101;
12'd1086 : tab2 = 23'b00001110011001110101010;
12'd1087 : tab2 = 23'b00001110010001100011101;
12'd1088 : tab2 = 23'b00001110001001010010001;
12'd1089 : tab2 = 23'b00001110000001000000111;
12'd1090 : tab2 = 23'b00001101111000110000101;
12'd1091 : tab2 = 23'b00001101110000100000100;
12'd1092 : tab2 = 23'b00001101101000010000101;
12'd1093 : tab2 = 23'b00001101100000000001010;
12'd1094 : tab2 = 23'b00001101010111110010110;
12'd1095 : tab2 = 23'b00001101001111100100000;
12'd1096 : tab2 = 23'b00001101000111010110000;
12'd1097 : tab2 = 23'b00001100111111001000100;
12'd1098 : tab2 = 23'b00001100110110111011011;
12'd1099 : tab2 = 23'b00001100101110101110100;
12'd1100 : tab2 = 23'b00001100100110100010001;
12'd1101 : tab2 = 23'b00001100011110010110010;
12'd1102 : tab2 = 23'b00001100010110001010111;
12'd1103 : tab2 = 23'b00001100001101111111100;
12'd1104 : tab2 = 23'b00001100000101110100110;
12'd1105 : tab2 = 23'b00001011111101101010101;
12'd1106 : tab2 = 23'b00001011110101100000101;
12'd1107 : tab2 = 23'b00001011101101010111011;
12'd1108 : tab2 = 23'b00001011100101001110010;
12'd1109 : tab2 = 23'b00001011011101000101101;
12'd1110 : tab2 = 23'b00001011010100111101001;
12'd1111 : tab2 = 23'b00001011001100110101011;
12'd1112 : tab2 = 23'b00001011000100101110010;
12'd1113 : tab2 = 23'b00001010111100100111010;
12'd1114 : tab2 = 23'b00001010110100100000100;
12'd1115 : tab2 = 23'b00001010101100011010011;
12'd1116 : tab2 = 23'b00001010100100010100101;
12'd1117 : tab2 = 23'b00001010011100001111100;
12'd1118 : tab2 = 23'b00001010010100001010011;
12'd1119 : tab2 = 23'b00001010001100000101110;
12'd1120 : tab2 = 23'b00001010000100000001111;
12'd1121 : tab2 = 23'b00001001111011111110010;
12'd1122 : tab2 = 23'b00001001110011111010101;
12'd1123 : tab2 = 23'b00001001101011110111110;
12'd1124 : tab2 = 23'b00001001100011110101010;
12'd1125 : tab2 = 23'b00001001011011110011011;
12'd1126 : tab2 = 23'b00001001010011110001011;
12'd1127 : tab2 = 23'b00001001001011110000001;
12'd1128 : tab2 = 23'b00001001000011101111100;
12'd1129 : tab2 = 23'b00001000111011101110110;
12'd1130 : tab2 = 23'b00001000110011101110110;
12'd1131 : tab2 = 23'b00001000101011101111000;
12'd1132 : tab2 = 23'b00001000100011101111110;
12'd1133 : tab2 = 23'b00001000011011110001001;
12'd1134 : tab2 = 23'b00001000010011110010011;
12'd1135 : tab2 = 23'b00001000001011110100100;
12'd1136 : tab2 = 23'b00001000000011110110101;
12'd1137 : tab2 = 23'b00000111111011111001101;
12'd1138 : tab2 = 23'b00000111110011111100100;
12'd1139 : tab2 = 23'b00000111101100000000011;
12'd1140 : tab2 = 23'b00000111100100000100000;
12'd1141 : tab2 = 23'b00000111011100001000101;
12'd1142 : tab2 = 23'b00000111010100001101001;
12'd1143 : tab2 = 23'b00000111001100010010010;
12'd1144 : tab2 = 23'b00000111000100010111110;
12'd1145 : tab2 = 23'b00000110111100011101110;
12'd1146 : tab2 = 23'b00000110110100100100000;
12'd1147 : tab2 = 23'b00000110101100101010110;
12'd1148 : tab2 = 23'b00000110100100110010001;
12'd1149 : tab2 = 23'b00000110011100111001011;
12'd1150 : tab2 = 23'b00000110010101000001010;
12'd1151 : tab2 = 23'b00000110001101001001101;
12'd1152 : tab2 = 23'b00000110000101010010001;
12'd1153 : tab2 = 23'b00000101111101011011010;
12'd1154 : tab2 = 23'b00000101110101100101000;
12'd1155 : tab2 = 23'b00000101101101101110111;
12'd1156 : tab2 = 23'b00000101100101111001000;
12'd1157 : tab2 = 23'b00000101011110000011101;
12'd1158 : tab2 = 23'b00000101010110001110100;
12'd1159 : tab2 = 23'b00000101001110011010001;
12'd1160 : tab2 = 23'b00000101000110100101110;
12'd1161 : tab2 = 23'b00000100111110110010000;
12'd1162 : tab2 = 23'b00000100110110111110101;
12'd1163 : tab2 = 23'b00000100101111001011100;
12'd1164 : tab2 = 23'b00000100100111011001010;
12'd1165 : tab2 = 23'b00000100011111100110100;
12'd1166 : tab2 = 23'b00000100010111110100111;
12'd1167 : tab2 = 23'b00000100010000000011110;
12'd1168 : tab2 = 23'b00000100001000010010010;
12'd1169 : tab2 = 23'b00000100000000100010000;
12'd1170 : tab2 = 23'b00000011111000110001011;
12'd1171 : tab2 = 23'b00000011110001000001011;
12'd1172 : tab2 = 23'b00000011101001010001101;
12'd1173 : tab2 = 23'b00000011100001100010110;
12'd1174 : tab2 = 23'b00000011011001110100001;
12'd1175 : tab2 = 23'b00000011010010000101101;
12'd1176 : tab2 = 23'b00000011001010010111101;
12'd1177 : tab2 = 23'b00000011000010101010010;
12'd1178 : tab2 = 23'b00000010111010111100111;
12'd1179 : tab2 = 23'b00000010110011001111110;
12'd1180 : tab2 = 23'b00000010101011100011010;
12'd1181 : tab2 = 23'b00000010100011110111011;
12'd1182 : tab2 = 23'b00000010011100001011110;
12'd1183 : tab2 = 23'b00000010010100100000011;
12'd1184 : tab2 = 23'b00000010001100110101100;
12'd1185 : tab2 = 23'b00000010000101001010101;
12'd1186 : tab2 = 23'b00000001111101100000100;
12'd1187 : tab2 = 23'b00000001110101110110110;
12'd1188 : tab2 = 23'b00000001101110001101011;
12'd1189 : tab2 = 23'b00000001100110100100001;
12'd1190 : tab2 = 23'b00000001011110111011101;
12'd1191 : tab2 = 23'b00000001010111010011011;
12'd1192 : tab2 = 23'b00000001001111101011100;
12'd1193 : tab2 = 23'b00000001001000000011111;
12'd1194 : tab2 = 23'b00000001000000011100101;
12'd1195 : tab2 = 23'b00000000111000110101111;
12'd1196 : tab2 = 23'b00000000110001001111101;
12'd1197 : tab2 = 23'b00000000101001101001010;
12'd1198 : tab2 = 23'b00000000100010000011110;
12'd1199 : tab2 = 23'b00000000011010011110100;
12'd1200 : tab2 = 23'b00000000010010111001110;
12'd1201 : tab2 = 23'b00000000001011010100111;
12'd1202 : tab2 = 23'b00000000000011110000101;
12'd1203 : tab2 = 23'b11111111111000011001110;
12'd1204 : tab2 = 23'b11111111101001010011100;
12'd1205 : tab2 = 23'b11111111011010001100110;
12'd1206 : tab2 = 23'b11111111001011000111101;
12'd1207 : tab2 = 23'b11111110111100000011000;
12'd1208 : tab2 = 23'b11111110101100111110110;
12'd1209 : tab2 = 23'b11111110011101111011101;
12'd1210 : tab2 = 23'b11111110001110111001000;
12'd1211 : tab2 = 23'b11111101111111110111100;
12'd1212 : tab2 = 23'b11111101110000110111010;
12'd1213 : tab2 = 23'b11111101100001110110011;
12'd1214 : tab2 = 23'b11111101010010110110110;
12'd1215 : tab2 = 23'b11111101000011111000010;
12'd1216 : tab2 = 23'b11111100110100111010010;
12'd1217 : tab2 = 23'b11111100100101111101000;
12'd1218 : tab2 = 23'b11111100010111000000000;
12'd1219 : tab2 = 23'b11111100001000000100100;
12'd1220 : tab2 = 23'b11111011111001001001100;
12'd1221 : tab2 = 23'b11111011101010001111010;
12'd1222 : tab2 = 23'b11111011011011010101001;
12'd1223 : tab2 = 23'b11111011001100011100111;
12'd1224 : tab2 = 23'b11111010111101100100111;
12'd1225 : tab2 = 23'b11111010101110101101000;
12'd1226 : tab2 = 23'b11111010011111110110100;
12'd1227 : tab2 = 23'b11111010010001000000011;
12'd1228 : tab2 = 23'b11111010000010001011100;
12'd1229 : tab2 = 23'b11111001110011010110101;
12'd1230 : tab2 = 23'b11111001100100100010101;
12'd1231 : tab2 = 23'b11111001010101110000000;
12'd1232 : tab2 = 23'b11111001000110111101010;
12'd1233 : tab2 = 23'b11111000111000001011100;
12'd1234 : tab2 = 23'b11111000101001011011000;
12'd1235 : tab2 = 23'b11111000011010101010000;
12'd1236 : tab2 = 23'b11111000001011111011000;
12'd1237 : tab2 = 23'b11110111111101001100011;
12'd1238 : tab2 = 23'b11110111101110011110001;
12'd1239 : tab2 = 23'b11110111011111110000111;
12'd1240 : tab2 = 23'b11110111010001000100000;
12'd1241 : tab2 = 23'b11110111000010011000100;
12'd1242 : tab2 = 23'b11110110110011101101001;
12'd1243 : tab2 = 23'b11110110100101000011000;
12'd1244 : tab2 = 23'b11110110010110011000010;
12'd1245 : tab2 = 23'b11110110000111101111101;
12'd1246 : tab2 = 23'b11110101111001000111010;
12'd1247 : tab2 = 23'b11110101101010011111110;
12'd1248 : tab2 = 23'b11110101011011111000110;
12'd1249 : tab2 = 23'b11110101001101010010110;
12'd1250 : tab2 = 23'b11110100111110101101011;
12'd1251 : tab2 = 23'b11110100110000001000010;
12'd1252 : tab2 = 23'b11110100100001100100100;
12'd1253 : tab2 = 23'b11110100010011000000111;
12'd1254 : tab2 = 23'b11110100000100011110010;
12'd1255 : tab2 = 23'b11110011110101111100001;
12'd1256 : tab2 = 23'b11110011100111011010110;
12'd1257 : tab2 = 23'b11110011011000111010010;
12'd1258 : tab2 = 23'b11110011001010011010011;
12'd1259 : tab2 = 23'b11110010111011111011110;
12'd1260 : tab2 = 23'b11110010101101011101000;
12'd1261 : tab2 = 23'b11110010011110111110111;
12'd1262 : tab2 = 23'b11110010010000100010001;
12'd1263 : tab2 = 23'b11110010000010000101111;
12'd1264 : tab2 = 23'b11110001110011101001101;
12'd1265 : tab2 = 23'b11110001100101001110100;
12'd1266 : tab2 = 23'b11110001010110110100001;
12'd1267 : tab2 = 23'b11110001001000011011000;
12'd1268 : tab2 = 23'b11110000111010000010011;
12'd1269 : tab2 = 23'b11110000101011101001101;
12'd1270 : tab2 = 23'b11110000011101010010011;
12'd1271 : tab2 = 23'b11110000001110111011101;
12'd1272 : tab2 = 23'b11110000000000100101010;
12'd1273 : tab2 = 23'b11101111110010001111101;
12'd1274 : tab2 = 23'b11101111100011111011010;
12'd1275 : tab2 = 23'b11101111010101100111001;
12'd1276 : tab2 = 23'b11101111000111010011110;
12'd1277 : tab2 = 23'b11101110111001000001100;
12'd1278 : tab2 = 23'b11101110101010101111000;
12'd1279 : tab2 = 23'b11101110011100011101111;
12'd1280 : tab2 = 23'b11101110001110001101100;
12'd1281 : tab2 = 23'b11101101111111111101110;
12'd1282 : tab2 = 23'b11101101110001101110001;
12'd1283 : tab2 = 23'b11101101100011011111100;
12'd1284 : tab2 = 23'b11101101010101010010001;
12'd1285 : tab2 = 23'b11101101000111000100010;
12'd1286 : tab2 = 23'b11101100111000111000001;
12'd1287 : tab2 = 23'b11101100101010101100000;
12'd1288 : tab2 = 23'b11101100011100100001000;
12'd1289 : tab2 = 23'b11101100001110010111000;
12'd1290 : tab2 = 23'b11101100000000001100101;
12'd1291 : tab2 = 23'b11101011110010000011110;
12'd1292 : tab2 = 23'b11101011100011111011000;
12'd1293 : tab2 = 23'b11101011010101110011010;
12'd1294 : tab2 = 23'b11101011000111101100101;
12'd1295 : tab2 = 23'b11101010111001100101110;
12'd1296 : tab2 = 23'b11101010101011100000000;
12'd1297 : tab2 = 23'b11101010011101011011001;
12'd1298 : tab2 = 23'b11101010001111010111000;
12'd1299 : tab2 = 23'b11101010000001010011000;
12'd1300 : tab2 = 23'b11101001110011001111111;
12'd1301 : tab2 = 23'b11101001100101001101111;
12'd1302 : tab2 = 23'b11101001010111001100001;
12'd1303 : tab2 = 23'b11101001001001001010100;
12'd1304 : tab2 = 23'b11101000111011001010001;
12'd1305 : tab2 = 23'b11101000101101001011000;
12'd1306 : tab2 = 23'b11101000011111001011110;
12'd1307 : tab2 = 23'b11101000010001001101101;
12'd1308 : tab2 = 23'b11101000000011001111111;
12'd1309 : tab2 = 23'b11100111110101010010110;
12'd1310 : tab2 = 23'b11100111100111010110001;
12'd1311 : tab2 = 23'b11100111011001011010100;
12'd1312 : tab2 = 23'b11100111001011011111101;
12'd1313 : tab2 = 23'b11100110111101100100111;
12'd1314 : tab2 = 23'b11100110101111101011011;
12'd1315 : tab2 = 23'b11100110100001110010101;
12'd1316 : tab2 = 23'b11100110010011111010000;
12'd1317 : tab2 = 23'b11100110000110000010001;
12'd1318 : tab2 = 23'b11100101111000001011000;
12'd1319 : tab2 = 23'b11100101101010010101001;
12'd1320 : tab2 = 23'b11100101011100011111000;
12'd1321 : tab2 = 23'b11100101001110101010000;
12'd1322 : tab2 = 23'b11100101000000110101011;
12'd1323 : tab2 = 23'b11100100110011000001111;
12'd1324 : tab2 = 23'b11100100100101001110001;
12'd1325 : tab2 = 23'b11100100010111011100001;
12'd1326 : tab2 = 23'b11100100001001101010010;
12'd1327 : tab2 = 23'b11100011111011111000110;
12'd1328 : tab2 = 23'b11100011101110001000010;
12'd1329 : tab2 = 23'b11100011100000011000101;
12'd1330 : tab2 = 23'b11100011010010101001011;
12'd1331 : tab2 = 23'b11100011000100111011000;
12'd1332 : tab2 = 23'b11100010110111001101001;
12'd1333 : tab2 = 23'b11100010101001011111011;
12'd1334 : tab2 = 23'b11100010011011110010110;
12'd1335 : tab2 = 23'b11100010001110000111000;
12'd1336 : tab2 = 23'b11100010000000011011111;
12'd1337 : tab2 = 23'b11100001110010110001011;
12'd1338 : tab2 = 23'b11100001100101000110110;
12'd1339 : tab2 = 23'b11100001010111011101011;
12'd1340 : tab2 = 23'b11100001001001110101001;
12'd1341 : tab2 = 23'b11100000111100001100101;
12'd1342 : tab2 = 23'b11100000101110100101011;
12'd1343 : tab2 = 23'b11100000100000111110111;
12'd1344 : tab2 = 23'b11100000010011011000100;
12'd1345 : tab2 = 23'b11100000000101110010010;
12'd1346 : tab2 = 23'b11011111111000001101111;
12'd1347 : tab2 = 23'b11011111101010101001101;
12'd1348 : tab2 = 23'b11011111011101000110001;
12'd1349 : tab2 = 23'b11011111001111100011000;
12'd1350 : tab2 = 23'b11011111000010000000111;
12'd1351 : tab2 = 23'b11011110110100011111000;
12'd1352 : tab2 = 23'b11011110100110111101111;
12'd1353 : tab2 = 23'b11011110011001011110000;
12'd1354 : tab2 = 23'b11011110001011111101110;
12'd1355 : tab2 = 23'b11011101111110011110110;
12'd1356 : tab2 = 23'b11011101110001000000000;
12'd1357 : tab2 = 23'b11011101100011100010010;
12'd1358 : tab2 = 23'b11011101010110000101000;
12'd1359 : tab2 = 23'b11011101001000100111110;
12'd1360 : tab2 = 23'b11011100111011001100011;
12'd1361 : tab2 = 23'b11011100101101110001010;
12'd1362 : tab2 = 23'b11011100100000010110010;
12'd1363 : tab2 = 23'b11011100010010111100011;
12'd1364 : tab2 = 23'b11011100000101100010110;
12'd1365 : tab2 = 23'b11011011111000001001100;
12'd1366 : tab2 = 23'b11011011101010110001101;
12'd1367 : tab2 = 23'b11011011011101011010001;
12'd1368 : tab2 = 23'b11011011010000000011000;
12'd1369 : tab2 = 23'b11011011000010101100100;
12'd1370 : tab2 = 23'b11011010110101010111001;
12'd1371 : tab2 = 23'b11011010101000000001100;
12'd1372 : tab2 = 23'b11011010011010101101000;
12'd1373 : tab2 = 23'b11011010001101011001011;
12'd1374 : tab2 = 23'b11011010000000000110010;
12'd1375 : tab2 = 23'b11011001110010110011111;
12'd1376 : tab2 = 23'b11011001100101100001011;
12'd1377 : tab2 = 23'b11011001011000010000011;
12'd1378 : tab2 = 23'b11011001001010111111010;
12'd1379 : tab2 = 23'b11011000111101101111010;
12'd1380 : tab2 = 23'b11011000110000100000000;
12'd1381 : tab2 = 23'b11011000100011010001011;
12'd1382 : tab2 = 23'b11011000010110000011000;
12'd1383 : tab2 = 23'b11011000001000110100110;
12'd1384 : tab2 = 23'b11010111111011100111110;
12'd1385 : tab2 = 23'b11010111101110011011101;
12'd1386 : tab2 = 23'b11010111100001001111100;
12'd1387 : tab2 = 23'b11010111010100000101010;
12'd1388 : tab2 = 23'b11010111000110111001111;
12'd1389 : tab2 = 23'b11010110111001110000001;
12'd1390 : tab2 = 23'b11010110101100100110110;
12'd1391 : tab2 = 23'b11010110011111011101110;
12'd1392 : tab2 = 23'b11010110010010010110011;
12'd1393 : tab2 = 23'b11010110000101001110010;
12'd1394 : tab2 = 23'b11010101111000000111011;
12'd1395 : tab2 = 23'b11010101101011000001000;
12'd1396 : tab2 = 23'b11010101011101111011100;
12'd1397 : tab2 = 23'b11010101010000110110001;
12'd1398 : tab2 = 23'b11010101000011110001100;
12'd1399 : tab2 = 23'b11010100110110101110011;
12'd1400 : tab2 = 23'b11010100101001101010101;
12'd1401 : tab2 = 23'b11010100011100101000001;
12'd1402 : tab2 = 23'b11010100001111100110010;
12'd1403 : tab2 = 23'b11010100000010100100100;
12'd1404 : tab2 = 23'b11010011110101100011100;
12'd1405 : tab2 = 23'b11010011101000100010111;
12'd1406 : tab2 = 23'b11010011011011100011110;
12'd1407 : tab2 = 23'b11010011001110100100111;
12'd1408 : tab2 = 23'b11010011000001100110101;
12'd1409 : tab2 = 23'b11010010110100101000101;
12'd1410 : tab2 = 23'b11010010100111101010111;
12'd1411 : tab2 = 23'b11010010011010101110001;
12'd1412 : tab2 = 23'b11010010001101110010011;
12'd1413 : tab2 = 23'b11010010000000110111001;
12'd1414 : tab2 = 23'b11010001110011111100001;
12'd1415 : tab2 = 23'b11010001100111000001110;
12'd1416 : tab2 = 23'b11010001011010001000001;
12'd1417 : tab2 = 23'b11010001001101001111000;
12'd1418 : tab2 = 23'b11010001000000010110011;
12'd1419 : tab2 = 23'b11010000110011011110111;
12'd1420 : tab2 = 23'b11010000100110100111100;
12'd1421 : tab2 = 23'b11010000011001110000110;
12'd1422 : tab2 = 23'b11010000001100111010010;
12'd1423 : tab2 = 23'b11010000000000000101000;
12'd1424 : tab2 = 23'b11001111110011001111111;
12'd1425 : tab2 = 23'b11001111100110011100000;
12'd1426 : tab2 = 23'b11001111011001101000010;
12'd1427 : tab2 = 23'b11001111001100110100101;
12'd1428 : tab2 = 23'b11001111000000000010010;
12'd1429 : tab2 = 23'b11001110110011010000101;
12'd1430 : tab2 = 23'b11001110100110011111001;
12'd1431 : tab2 = 23'b11001110011001101110011;
12'd1432 : tab2 = 23'b11001110001100111101111;
12'd1433 : tab2 = 23'b11001110000000001110011;
12'd1434 : tab2 = 23'b11001101110011011111101;
12'd1435 : tab2 = 23'b11001101100110110001000;
12'd1436 : tab2 = 23'b11001101011010000011011;
12'd1437 : tab2 = 23'b11001101001101010110001;
12'd1438 : tab2 = 23'b11001101000000101001010;
12'd1439 : tab2 = 23'b11001100110011111101101;
12'd1440 : tab2 = 23'b11001100100111010001101;
12'd1441 : tab2 = 23'b11001100011010100110110;
12'd1442 : tab2 = 23'b11001100001101111100100;
12'd1443 : tab2 = 23'b11001100000001010010100;
12'd1444 : tab2 = 23'b11001011110100101001001;
12'd1445 : tab2 = 23'b11001011101000000000111;
12'd1446 : tab2 = 23'b11001011011011011000100;
12'd1447 : tab2 = 23'b11001011001110110001001;
12'd1448 : tab2 = 23'b11001011000010001010011;
12'd1449 : tab2 = 23'b11001010110101100100000;
12'd1450 : tab2 = 23'b11001010101000111101111;
12'd1451 : tab2 = 23'b11001010011100011000110;
12'd1452 : tab2 = 23'b11001010001111110100111;
12'd1453 : tab2 = 23'b11001010000011010000001;
12'd1454 : tab2 = 23'b11001001110110101100101;
12'd1455 : tab2 = 23'b11001001101010001010010;
12'd1456 : tab2 = 23'b11001001011101101000001;
12'd1457 : tab2 = 23'b11001001010001000110000;
12'd1458 : tab2 = 23'b11001001000100100100110;
12'd1459 : tab2 = 23'b11001000111000000100101;
12'd1460 : tab2 = 23'b11001000101011100100101;
12'd1461 : tab2 = 23'b11001000011111000100110;
12'd1462 : tab2 = 23'b11001000010010100101111;
12'd1463 : tab2 = 23'b11001000000110000111111;
12'd1464 : tab2 = 23'b11000111111001101010001;
12'd1465 : tab2 = 23'b11000111101101001100100;
12'd1466 : tab2 = 23'b11000111100000110000010;
12'd1467 : tab2 = 23'b11000111010100010100000;
12'd1468 : tab2 = 23'b11000111000111111000111;
12'd1469 : tab2 = 23'b11000110111011011110000;
12'd1470 : tab2 = 23'b11000110101111000011011;
12'd1471 : tab2 = 23'b11000110100010101001110;
12'd1472 : tab2 = 23'b11000110010110010000101;
12'd1473 : tab2 = 23'b11000110001001110111111;
12'd1474 : tab2 = 23'b11000101111101011111100;
12'd1475 : tab2 = 23'b11000101110001001000101;
12'd1476 : tab2 = 23'b11000101100100110001000;
12'd1477 : tab2 = 23'b11000101011000011010101;
12'd1478 : tab2 = 23'b11000101001100000100110;
12'd1479 : tab2 = 23'b11000100111111101111010;
12'd1480 : tab2 = 23'b11000100110011011011010;
12'd1481 : tab2 = 23'b11000100100111000110100;
12'd1482 : tab2 = 23'b11000100011010110011000;
12'd1483 : tab2 = 23'b11000100001110100000100;
12'd1484 : tab2 = 23'b11000100000010001101011;
12'd1485 : tab2 = 23'b11000011110101111011110;
12'd1486 : tab2 = 23'b11000011101001101010011;
12'd1487 : tab2 = 23'b11000011011101011001110;
12'd1488 : tab2 = 23'b11000011010001001001001;
12'd1489 : tab2 = 23'b11000011000100111001101;
12'd1490 : tab2 = 23'b11000010111000101010100;
12'd1491 : tab2 = 23'b11000010101100011011101;
12'd1492 : tab2 = 23'b11000010100000001101101;
12'd1493 : tab2 = 23'b11000010010100000000001;
12'd1494 : tab2 = 23'b11000010000111110011001;
12'd1495 : tab2 = 23'b11000001111011100111000;
12'd1496 : tab2 = 23'b11000001101111011010111;
12'd1497 : tab2 = 23'b11000001100011001111100;
12'd1498 : tab2 = 23'b11000001010111000101000;
12'd1499 : tab2 = 23'b11000001001010111010110;
12'd1500 : tab2 = 23'b11000000111110110001000;
12'd1501 : tab2 = 23'b11000000110010101000001;
12'd1502 : tab2 = 23'b11000000100110011111011;
12'd1503 : tab2 = 23'b11000000011010010111011;
12'd1504 : tab2 = 23'b11000000001110010000000;
12'd1505 : tab2 = 23'b11000000000010001001000;
12'd1506 : tab2 = 23'b10111111110110000010011;
12'd1507 : tab2 = 23'b10111111101001111101001;
12'd1508 : tab2 = 23'b10111111011101110111111;
12'd1509 : tab2 = 23'b10111111010001110010110;
12'd1510 : tab2 = 23'b10111111000101101110101;
12'd1511 : tab2 = 23'b10111110111001101011011;
12'd1512 : tab2 = 23'b10111110101101100111110;
12'd1513 : tab2 = 23'b10111110100001100101011;
12'd1514 : tab2 = 23'b10111110010101100011011;
12'd1515 : tab2 = 23'b10111110001001100001011;
12'd1516 : tab2 = 23'b10111101111101100000100;
12'd1517 : tab2 = 23'b10111101110001100000010;
12'd1518 : tab2 = 23'b10111101100101100000011;
12'd1519 : tab2 = 23'b10111101011001100000111;
12'd1520 : tab2 = 23'b10111101001101100010101;
12'd1521 : tab2 = 23'b10111101000001100011110;
12'd1522 : tab2 = 23'b10111100110101100101111;
12'd1523 : tab2 = 23'b10111100101001101001001;
12'd1524 : tab2 = 23'b10111100011101101100100;
12'd1525 : tab2 = 23'b10111100010001110000010;
12'd1526 : tab2 = 23'b10111100000101110100100;
12'd1527 : tab2 = 23'b10111011111001111001111;
12'd1528 : tab2 = 23'b10111011101101111111001;
12'd1529 : tab2 = 23'b10111011100010000101010;
12'd1530 : tab2 = 23'b10111011010110001011110;
12'd1531 : tab2 = 23'b10111011001010010010011;
12'd1532 : tab2 = 23'b10111010111110011010001;
12'd1533 : tab2 = 23'b10111010110010100010100;
12'd1534 : tab2 = 23'b10111010100110101011001;
12'd1535 : tab2 = 23'b10111010011010110100010;
12'd1536 : tab2 = 23'b10111010001110111110100;
12'd1537 : tab2 = 23'b10111010000011001000010;
12'd1538 : tab2 = 23'b10111001110111010010110;
12'd1539 : tab2 = 23'b10111001101011011110010;
12'd1540 : tab2 = 23'b10111001011111101010010;
12'd1541 : tab2 = 23'b10111001010011110110111;
12'd1542 : tab2 = 23'b10111001001000000011001;
12'd1543 : tab2 = 23'b10111000111100010000110;
12'd1544 : tab2 = 23'b10111000110000011110111;
12'd1545 : tab2 = 23'b10111000100100101101010;
12'd1546 : tab2 = 23'b10111000011000111100000;
12'd1547 : tab2 = 23'b10111000001101001011110;
12'd1548 : tab2 = 23'b10111000000001011100000;
12'd1549 : tab2 = 23'b10110111110101101100100;
12'd1550 : tab2 = 23'b10110111101001111101011;
12'd1551 : tab2 = 23'b10110111011110001111001;
12'd1552 : tab2 = 23'b10110111010010100001000;
12'd1553 : tab2 = 23'b10110111000110110011101;
12'd1554 : tab2 = 23'b10110110111011000111001;
12'd1555 : tab2 = 23'b10110110101111011010110;
12'd1556 : tab2 = 23'b10110110100011101111001;
12'd1557 : tab2 = 23'b10110110011000000011110;
12'd1558 : tab2 = 23'b10110110001100011001001;
12'd1559 : tab2 = 23'b10110110000000101110100;
12'd1560 : tab2 = 23'b10110101110101000100101;
12'd1561 : tab2 = 23'b10110101101001011011100;
12'd1562 : tab2 = 23'b10110101011101110011010;
12'd1563 : tab2 = 23'b10110101010010001011000;
12'd1564 : tab2 = 23'b10110101000110100011010;
12'd1565 : tab2 = 23'b10110100111010111100100;
12'd1566 : tab2 = 23'b10110100101111010101100;
12'd1567 : tab2 = 23'b10110100100011101111101;
12'd1568 : tab2 = 23'b10110100011000001001100;
12'd1569 : tab2 = 23'b10110100001100100100100;
12'd1570 : tab2 = 23'b10110100000001000000001;
12'd1571 : tab2 = 23'b10110011110101011011111;
12'd1572 : tab2 = 23'b10110011101001111000011;
12'd1573 : tab2 = 23'b10110011011110010101011;
12'd1574 : tab2 = 23'b10110011010010110010101;
12'd1575 : tab2 = 23'b10110011000111010000100;
12'd1576 : tab2 = 23'b10110010111011101111001;
12'd1577 : tab2 = 23'b10110010110000001101110;
12'd1578 : tab2 = 23'b10110010100100101101101;
12'd1579 : tab2 = 23'b10110010011001001101100;
12'd1580 : tab2 = 23'b10110010001101101110001;
12'd1581 : tab2 = 23'b10110010000010001111100;
12'd1582 : tab2 = 23'b10110001110110110000011;
12'd1583 : tab2 = 23'b10110001101011010010111;
12'd1584 : tab2 = 23'b10110001011111110101101;
12'd1585 : tab2 = 23'b10110001010100011000100;
12'd1586 : tab2 = 23'b10110001001000111100000;
12'd1587 : tab2 = 23'b10110000111101011111101;
12'd1588 : tab2 = 23'b10110000110010000100011;
12'd1589 : tab2 = 23'b10110000100110101001011;
12'd1590 : tab2 = 23'b10110000011011001110111;
12'd1591 : tab2 = 23'b10110000001111110101001;
12'd1592 : tab2 = 23'b10110000000100011011100;
12'd1593 : tab2 = 23'b10101111111001000010100;
12'd1594 : tab2 = 23'b10101111101101101010100;
12'd1595 : tab2 = 23'b10101111100010010010000;
12'd1596 : tab2 = 23'b10101111010110111011010;
12'd1597 : tab2 = 23'b10101111001011100100000;
12'd1598 : tab2 = 23'b10101111000000001101110;
12'd1599 : tab2 = 23'b10101110110100110111101;
12'd1600 : tab2 = 23'b10101110101001100010001;
12'd1601 : tab2 = 23'b10101110011110001101011;
12'd1602 : tab2 = 23'b10101110010010111000101;
12'd1603 : tab2 = 23'b10101110000111100100101;
12'd1604 : tab2 = 23'b10101101111100010001010;
12'd1605 : tab2 = 23'b10101101110000111101111;
12'd1606 : tab2 = 23'b10101101100101101011111;
12'd1607 : tab2 = 23'b10101101011010011001111;
12'd1608 : tab2 = 23'b10101101001111001000000;
12'd1609 : tab2 = 23'b10101101000011110111010;
12'd1610 : tab2 = 23'b10101100111000100110110;
12'd1611 : tab2 = 23'b10101100101101010110011;
12'd1612 : tab2 = 23'b10101100100010000111000;
12'd1613 : tab2 = 23'b10101100010110110111111;
12'd1614 : tab2 = 23'b10101100001011101001110;
12'd1615 : tab2 = 23'b10101100000000011011101;
12'd1616 : tab2 = 23'b10101011110101001110010;
12'd1617 : tab2 = 23'b10101011101010000000110;
12'd1618 : tab2 = 23'b10101011011110110100011;
12'd1619 : tab2 = 23'b10101011010011101000001;
12'd1620 : tab2 = 23'b10101011001000011100110;
12'd1621 : tab2 = 23'b10101010111101010001110;
12'd1622 : tab2 = 23'b10101010110010000110111;
12'd1623 : tab2 = 23'b10101010100110111101001;
12'd1624 : tab2 = 23'b10101010011011110011000;
12'd1625 : tab2 = 23'b10101010010000101010001;
12'd1626 : tab2 = 23'b10101010000101100001101;
12'd1627 : tab2 = 23'b10101001111010011001000;
12'd1628 : tab2 = 23'b10101001101111010001011;
12'd1629 : tab2 = 23'b10101001100100001010011;
12'd1630 : tab2 = 23'b10101001011001000011001;
12'd1631 : tab2 = 23'b10101001001101111101000;
12'd1632 : tab2 = 23'b10101001000010110111100;
12'd1633 : tab2 = 23'b10101000110111110010001;
12'd1634 : tab2 = 23'b10101000101100101101010;
12'd1635 : tab2 = 23'b10101000100001101001010;
12'd1636 : tab2 = 23'b10101000010110100101010;
12'd1637 : tab2 = 23'b10101000001011100001111;
12'd1638 : tab2 = 23'b10101000000000011110110;
12'd1639 : tab2 = 23'b10100111110101011100100;
12'd1640 : tab2 = 23'b10100111101010011010010;
12'd1641 : tab2 = 23'b10100111011111011000111;
12'd1642 : tab2 = 23'b10100111010100010111110;
12'd1643 : tab2 = 23'b10100111001001010111110;
12'd1644 : tab2 = 23'b10100110111110010111011;
12'd1645 : tab2 = 23'b10100110110011010111111;
12'd1646 : tab2 = 23'b10100110101000011000111;
12'd1647 : tab2 = 23'b10100110011101011001111;
12'd1648 : tab2 = 23'b10100110010010011100011;
12'd1649 : tab2 = 23'b10100110000111011110001;
12'd1650 : tab2 = 23'b10100101111100100001001;
12'd1651 : tab2 = 23'b10100101110001100100100;
12'd1652 : tab2 = 23'b10100101100110101000010;
12'd1653 : tab2 = 23'b10100101011011101100100;
12'd1654 : tab2 = 23'b10100101010000110001000;
12'd1655 : tab2 = 23'b10100101000101110110100;
12'd1656 : tab2 = 23'b10100100111010111100001;
12'd1657 : tab2 = 23'b10100100110000000010000;
12'd1658 : tab2 = 23'b10100100100101001000111;
12'd1659 : tab2 = 23'b10100100011010001111111;
12'd1660 : tab2 = 23'b10100100001111010111101;
12'd1661 : tab2 = 23'b10100100000100011111100;
12'd1662 : tab2 = 23'b10100011111001100111111;
12'd1663 : tab2 = 23'b10100011101110110000100;
12'd1664 : tab2 = 23'b10100011100011111010001;
12'd1665 : tab2 = 23'b10100011011001000100000;
12'd1666 : tab2 = 23'b10100011001110001110011;
12'd1667 : tab2 = 23'b10100011000011011001001;
12'd1668 : tab2 = 23'b10100010111000100100110;
12'd1669 : tab2 = 23'b10100010101101110000100;
12'd1670 : tab2 = 23'b10100010100010111100100;
12'd1671 : tab2 = 23'b10100010011000001001010;
12'd1672 : tab2 = 23'b10100010001101010110011;
12'd1673 : tab2 = 23'b10100010000010100011111;
12'd1674 : tab2 = 23'b10100001110111110010010;
12'd1675 : tab2 = 23'b10100001101101000000011;
12'd1676 : tab2 = 23'b10100001100010001111101;
12'd1677 : tab2 = 23'b10100001010111011111000;
12'd1678 : tab2 = 23'b10100001001100101110111;
12'd1679 : tab2 = 23'b10100001000001111111100;
12'd1680 : tab2 = 23'b10100000110111010000011;
12'd1681 : tab2 = 23'b10100000101100100001101;
12'd1682 : tab2 = 23'b10100000100001110011001;
12'd1683 : tab2 = 23'b10100000010111000101101;
12'd1684 : tab2 = 23'b10100000001100011000000;
12'd1685 : tab2 = 23'b10100000000001101011011;
12'd1686 : tab2 = 23'b10011111110110111110110;
12'd1687 : tab2 = 23'b10011111101100010010111;
12'd1688 : tab2 = 23'b10011111100001100111010;
12'd1689 : tab2 = 23'b10011111010110111100101;
12'd1690 : tab2 = 23'b10011111001100010010000;
12'd1691 : tab2 = 23'b10011111000001100111101;
12'd1692 : tab2 = 23'b10011110110110111110011;
12'd1693 : tab2 = 23'b10011110101100010100101;
12'd1694 : tab2 = 23'b10011110100001101100001;
12'd1695 : tab2 = 23'b10011110010111000011110;
12'd1696 : tab2 = 23'b10011110001100011011111;
12'd1697 : tab2 = 23'b10011110000001110100110;
12'd1698 : tab2 = 23'b10011101110111001101110;
12'd1699 : tab2 = 23'b10011101101100100111010;
12'd1700 : tab2 = 23'b10011101100010000001100;
12'd1701 : tab2 = 23'b10011101010111011011111;
12'd1702 : tab2 = 23'b10011101001100110110010;
12'd1703 : tab2 = 23'b10011101000010010001111;
12'd1704 : tab2 = 23'b10011100110111101101101;
12'd1705 : tab2 = 23'b10011100101101001001111;
12'd1706 : tab2 = 23'b10011100100010100110011;
12'd1707 : tab2 = 23'b10011100011000000011100;
12'd1708 : tab2 = 23'b10011100001101100001100;
12'd1709 : tab2 = 23'b10011100000010111110110;
12'd1710 : tab2 = 23'b10011011111000011101110;
12'd1711 : tab2 = 23'b10011011101101111100101;
12'd1712 : tab2 = 23'b10011011100011011011111;
12'd1713 : tab2 = 23'b10011011011000111100000;
12'd1714 : tab2 = 23'b10011011001110011011111;
12'd1715 : tab2 = 23'b10011011000011111101000;
12'd1716 : tab2 = 23'b10011010111001011110000;
12'd1717 : tab2 = 23'b10011010101110111111010;
12'd1718 : tab2 = 23'b10011010100100100001110;
12'd1719 : tab2 = 23'b10011010011010000100001;
12'd1720 : tab2 = 23'b10011010001111100110110;
12'd1721 : tab2 = 23'b10011010000101001010011;
12'd1722 : tab2 = 23'b10011001111010101110010;
12'd1723 : tab2 = 23'b10011001110000010010010;
12'd1724 : tab2 = 23'b10011001100101110111010;
12'd1725 : tab2 = 23'b10011001011011011100011;
12'd1726 : tab2 = 23'b10011001010001000001110;
12'd1727 : tab2 = 23'b10011001000110100111101;
12'd1728 : tab2 = 23'b10011000111100001110100;
12'd1729 : tab2 = 23'b10011000110001110101010;
12'd1730 : tab2 = 23'b10011000100111011101000;
12'd1731 : tab2 = 23'b10011000011101000100110;
12'd1732 : tab2 = 23'b10011000010010101100110;
12'd1733 : tab2 = 23'b10011000001000010101000;
12'd1734 : tab2 = 23'b10010111111101111110001;
12'd1735 : tab2 = 23'b10010111110011101000011;
12'd1736 : tab2 = 23'b10010111101001010001111;
12'd1737 : tab2 = 23'b10010111011110111100011;
12'd1738 : tab2 = 23'b10010111010100100111001;
12'd1739 : tab2 = 23'b10010111001010010010110;
12'd1740 : tab2 = 23'b10010110111111111110101;
12'd1741 : tab2 = 23'b10010110110101101010101;
12'd1742 : tab2 = 23'b10010110101011010111000;
12'd1743 : tab2 = 23'b10010110100001000100001;
12'd1744 : tab2 = 23'b10010110010110110001100;
12'd1745 : tab2 = 23'b10010110001100011111100;
12'd1746 : tab2 = 23'b10010110000010001101111;
12'd1747 : tab2 = 23'b10010101110111111101001;
12'd1748 : tab2 = 23'b10010101101101101011111;
12'd1749 : tab2 = 23'b10010101100011011011111;
12'd1750 : tab2 = 23'b10010101011001001011110;
12'd1751 : tab2 = 23'b10010101001110111100001;
12'd1752 : tab2 = 23'b10010101000100101101001;
12'd1753 : tab2 = 23'b10010100111010011110101;
12'd1754 : tab2 = 23'b10010100110000010000001;
12'd1755 : tab2 = 23'b10010100100110000010100;
12'd1756 : tab2 = 23'b10010100011011110101010;
12'd1757 : tab2 = 23'b10010100010001101000001;
12'd1758 : tab2 = 23'b10010100000111011100000;
12'd1759 : tab2 = 23'b10010011111101001111100;
12'd1760 : tab2 = 23'b10010011110011000100001;
12'd1761 : tab2 = 23'b10010011101000111000011;
12'd1762 : tab2 = 23'b10010011011110101101101;
12'd1763 : tab2 = 23'b10010011010100100011110;
12'd1764 : tab2 = 23'b10010011001010011001101;
12'd1765 : tab2 = 23'b10010011000000010000010;
12'd1766 : tab2 = 23'b10010010110110000111001;
12'd1767 : tab2 = 23'b10010010101011111110100;
12'd1768 : tab2 = 23'b10010010100001110110001;
12'd1769 : tab2 = 23'b10010010010111101110001;
12'd1770 : tab2 = 23'b10010010001101100111011;
12'd1771 : tab2 = 23'b10010010000011100000001;
12'd1772 : tab2 = 23'b10010001111001011001001;
12'd1773 : tab2 = 23'b10010001101111010011100;
12'd1774 : tab2 = 23'b10010001100101001101110;
12'd1775 : tab2 = 23'b10010001011011001000100;
12'd1776 : tab2 = 23'b10010001010001000011110;
12'd1777 : tab2 = 23'b10010001000110111111011;
12'd1778 : tab2 = 23'b10010000111100111011011;
12'd1779 : tab2 = 23'b10010000110010110111101;
12'd1780 : tab2 = 23'b10010000101000110100011;
12'd1781 : tab2 = 23'b10010000011110110001110;
12'd1782 : tab2 = 23'b10010000010100101111101;
12'd1783 : tab2 = 23'b10010000001010101101110;
12'd1784 : tab2 = 23'b10010000000000101100000;
12'd1785 : tab2 = 23'b10001111110110101011001;
12'd1786 : tab2 = 23'b10001111101100101010010;
12'd1787 : tab2 = 23'b10001111100010101010001;
12'd1788 : tab2 = 23'b10001111011000101010011;
12'd1789 : tab2 = 23'b10001111001110101010101;
12'd1790 : tab2 = 23'b10001111000100101011111;
12'd1791 : tab2 = 23'b10001110111010101101011;
12'd1792 : tab2 = 23'b10001110110000101111000;
12'd1793 : tab2 = 23'b10001110100110110001100;
12'd1794 : tab2 = 23'b10001110011100110100001;
12'd1795 : tab2 = 23'b10001110010010110111001;
12'd1796 : tab2 = 23'b10001110001000111011000;
12'd1797 : tab2 = 23'b10001101111110111111000;
12'd1798 : tab2 = 23'b10001101110101000011010;
12'd1799 : tab2 = 23'b10001101101011000111111;
12'd1800 : tab2 = 23'b10001101100001001100111;
12'd1801 : tab2 = 23'b10001101010111010010011;
12'd1802 : tab2 = 23'b10001101001101011000111;
12'd1803 : tab2 = 23'b10001101000011011111000;
12'd1804 : tab2 = 23'b10001100111001100110010;
12'd1805 : tab2 = 23'b10001100101111101101001;
12'd1806 : tab2 = 23'b10001100100101110100100;
12'd1807 : tab2 = 23'b10001100011011111100101;
12'd1808 : tab2 = 23'b10001100010010000101010;
12'd1809 : tab2 = 23'b10001100001000001101110;
12'd1810 : tab2 = 23'b10001011111110010111001;
12'd1811 : tab2 = 23'b10001011110100100001000;
12'd1812 : tab2 = 23'b10001011101010101011001;
12'd1813 : tab2 = 23'b10001011100000110101110;
12'd1814 : tab2 = 23'b10001011010111000000101;
12'd1815 : tab2 = 23'b10001011001101001011100;
12'd1816 : tab2 = 23'b10001011000011010111011;
12'd1817 : tab2 = 23'b10001010111001100011100;
12'd1818 : tab2 = 23'b10001010101111110000010;
12'd1819 : tab2 = 23'b10001010100101111101011;
12'd1820 : tab2 = 23'b10001010011100001010011;
12'd1821 : tab2 = 23'b10001010010010011000010;
12'd1822 : tab2 = 23'b10001010001000100110011;
12'd1823 : tab2 = 23'b10001001111110110101000;
12'd1824 : tab2 = 23'b10001001110101000011111;
12'd1825 : tab2 = 23'b10001001101011010011101;
12'd1826 : tab2 = 23'b10001001100001100010110;
12'd1827 : tab2 = 23'b10001001010111110011010;
12'd1828 : tab2 = 23'b10001001001110000011111;
12'd1829 : tab2 = 23'b10001001000100010100101;
12'd1830 : tab2 = 23'b10001000111010100110011;
12'd1831 : tab2 = 23'b10001000110000111000000;
12'd1832 : tab2 = 23'b10001000100111001010011;
12'd1833 : tab2 = 23'b10001000011101011100101;
12'd1834 : tab2 = 23'b10001000010011101111111;
12'd1835 : tab2 = 23'b10001000001010000011010;
12'd1836 : tab2 = 23'b10001000000000010110110;
12'd1837 : tab2 = 23'b10000111110110101010110;
12'd1838 : tab2 = 23'b10000111101100111111011;
12'd1839 : tab2 = 23'b10000111100011010100101;
12'd1840 : tab2 = 23'b10000111011001101001100;
12'd1841 : tab2 = 23'b10000111001111111111110;
12'd1842 : tab2 = 23'b10000111000110010101111;
12'd1843 : tab2 = 23'b10000110111100101100110;
12'd1844 : tab2 = 23'b10000110110011000011010;
12'd1845 : tab2 = 23'b10000110101001011011000;
12'd1846 : tab2 = 23'b10000110011111110010011;
12'd1847 : tab2 = 23'b10000110010110001010010;
12'd1848 : tab2 = 23'b10000110001100100011000;
12'd1849 : tab2 = 23'b10000110000010111100001;
12'd1850 : tab2 = 23'b10000101111001010101010;
12'd1851 : tab2 = 23'b10000101101111101111010;
12'd1852 : tab2 = 23'b10000101100110001001001;
12'd1853 : tab2 = 23'b10000101011100100011011;
12'd1854 : tab2 = 23'b10000101010010111110110;
12'd1855 : tab2 = 23'b10000101001001011010001;
12'd1856 : tab2 = 23'b10000100111111110101111;
12'd1857 : tab2 = 23'b10000100110110010001111;
12'd1858 : tab2 = 23'b10000100101100101110011;
12'd1859 : tab2 = 23'b10000100100011001010111;
12'd1860 : tab2 = 23'b10000100011001101000101;
12'd1861 : tab2 = 23'b10000100010000000101111;
12'd1862 : tab2 = 23'b10000100000110100011111;
12'd1863 : tab2 = 23'b10000011111101000010011;
12'd1864 : tab2 = 23'b10000011110011100001100;
12'd1865 : tab2 = 23'b10000011101010000000001;
12'd1866 : tab2 = 23'b10000011100000100000000;
12'd1867 : tab2 = 23'b10000011010110111111111;
12'd1868 : tab2 = 23'b10000011001101100000101;
12'd1869 : tab2 = 23'b10000011000100000001010;
12'd1870 : tab2 = 23'b10000010111010100010000;
12'd1871 : tab2 = 23'b10000010110001000100000;
12'd1872 : tab2 = 23'b10000010100111100101100;
12'd1873 : tab2 = 23'b10000010011110000111110;
12'd1874 : tab2 = 23'b10000010010100101010101;
12'd1875 : tab2 = 23'b10000010001011001101111;
12'd1876 : tab2 = 23'b10000010000001110001100;
12'd1877 : tab2 = 23'b10000001111000010101001;
12'd1878 : tab2 = 23'b10000001101110111001001;
12'd1879 : tab2 = 23'b10000001100101011110000;
12'd1880 : tab2 = 23'b10000001011100000011000;
12'd1881 : tab2 = 23'b10000001010010101000001;
12'd1882 : tab2 = 23'b10000001001001001110011;
12'd1883 : tab2 = 23'b10000000111111110100101;
12'd1884 : tab2 = 23'b10000000110110011011000;
12'd1885 : tab2 = 23'b10000000101101000001100;
12'd1886 : tab2 = 23'b10000000100011101001000;
12'd1887 : tab2 = 23'b10000000011010010000110;
12'd1888 : tab2 = 23'b10000000010000111000110;
12'd1889 : tab2 = 23'b10000000000111100001001;
12'd1890 : tab2 = 23'b01111111111110001010001;
12'd1891 : tab2 = 23'b01111111110100110011001;
12'd1892 : tab2 = 23'b01111111101011011100101;
12'd1893 : tab2 = 23'b01111111100010000110011;
12'd1894 : tab2 = 23'b01111111011000110000110;
12'd1895 : tab2 = 23'b01111111001111011100000;
12'd1896 : tab2 = 23'b01111111000110000110111;
12'd1897 : tab2 = 23'b01111110111100110010100;
12'd1898 : tab2 = 23'b01111110110011011110100;
12'd1899 : tab2 = 23'b01111110101010001010011;
12'd1900 : tab2 = 23'b01111110100000110111001;
12'd1901 : tab2 = 23'b01111110010111100011111;
12'd1902 : tab2 = 23'b01111110001110010001110;
12'd1903 : tab2 = 23'b01111110000100111111000;
12'd1904 : tab2 = 23'b01111101111011101101001;
12'd1905 : tab2 = 23'b01111101110010011100001;
12'd1906 : tab2 = 23'b01111101101001001010100;
12'd1907 : tab2 = 23'b01111101011111111001111;
12'd1908 : tab2 = 23'b01111101010110101001011;
12'd1909 : tab2 = 23'b01111101001101011001111;
12'd1910 : tab2 = 23'b01111101000100001001101;
12'd1911 : tab2 = 23'b01111100111010111010011;
12'd1912 : tab2 = 23'b01111100110001101011100;
12'd1913 : tab2 = 23'b01111100101000011101000;
12'd1914 : tab2 = 23'b01111100011111001111000;
12'd1915 : tab2 = 23'b01111100010110000001000;
12'd1916 : tab2 = 23'b01111100001100110100000;
12'd1917 : tab2 = 23'b01111100000011100110111;
12'd1918 : tab2 = 23'b01111011111010011010101;
12'd1919 : tab2 = 23'b01111011110001001110001;
12'd1920 : tab2 = 23'b01111011101000000010000;
12'd1921 : tab2 = 23'b01111011011110110110100;
12'd1922 : tab2 = 23'b01111011010101101011010;
12'd1923 : tab2 = 23'b01111011001100100000100;
12'd1924 : tab2 = 23'b01111011000011010110010;
12'd1925 : tab2 = 23'b01111010111010001100001;
12'd1926 : tab2 = 23'b01111010110001000010001;
12'd1927 : tab2 = 23'b01111010100111111001001;
12'd1928 : tab2 = 23'b01111010011110110000001;
12'd1929 : tab2 = 23'b01111010010101100111001;
12'd1930 : tab2 = 23'b01111010001100011110111;
12'd1931 : tab2 = 23'b01111010000011010111001;
12'd1932 : tab2 = 23'b01111001111010001111101;
12'd1933 : tab2 = 23'b01111001110001001000010;
12'd1934 : tab2 = 23'b01111001101000000001110;
12'd1935 : tab2 = 23'b01111001011110111011101;
12'd1936 : tab2 = 23'b01111001010101110101100;
12'd1937 : tab2 = 23'b01111001001100101111011;
12'd1938 : tab2 = 23'b01111001000011101010010;
12'd1939 : tab2 = 23'b01111000111010100101010;
12'd1940 : tab2 = 23'b01111000110001100000111;
12'd1941 : tab2 = 23'b01111000101000011100101;
12'd1942 : tab2 = 23'b01111000011111011000111;
12'd1943 : tab2 = 23'b01111000010110010101010;
12'd1944 : tab2 = 23'b01111000001101010010001;
12'd1945 : tab2 = 23'b01111000000100001111001;
12'd1946 : tab2 = 23'b01110111111011001100110;
12'd1947 : tab2 = 23'b01110111110010001010101;
12'd1948 : tab2 = 23'b01110111101001001001001;
12'd1949 : tab2 = 23'b01110111100000001000000;
12'd1950 : tab2 = 23'b01110111010111000111000;
12'd1951 : tab2 = 23'b01110111001110000110100;
12'd1952 : tab2 = 23'b01110111000101000110011;
12'd1953 : tab2 = 23'b01110110111100000110101;
12'd1954 : tab2 = 23'b01110110110011000110111;
12'd1955 : tab2 = 23'b01110110101010000111101;
12'd1956 : tab2 = 23'b01110110100001001000111;
12'd1957 : tab2 = 23'b01110110011000001010100;
12'd1958 : tab2 = 23'b01110110001111001100100;
12'd1959 : tab2 = 23'b01110110000110001110101;
12'd1960 : tab2 = 23'b01110101111101010001011;
12'd1961 : tab2 = 23'b01110101110100010100010;
12'd1962 : tab2 = 23'b01110101101011010111111;
12'd1963 : tab2 = 23'b01110101100010011011100;
12'd1964 : tab2 = 23'b01110101011001011111100;
12'd1965 : tab2 = 23'b01110101010000100100000;
12'd1966 : tab2 = 23'b01110101000111101000101;
12'd1967 : tab2 = 23'b01110100111110101101111;
12'd1968 : tab2 = 23'b01110100110101110010110;
12'd1969 : tab2 = 23'b01110100101100111001000;
12'd1970 : tab2 = 23'b01110100100011111111100;
12'd1971 : tab2 = 23'b01110100011011000110001;
12'd1972 : tab2 = 23'b01110100010010001100110;
12'd1973 : tab2 = 23'b01110100001001010011111;
12'd1974 : tab2 = 23'b01110100000000011100000;
12'd1975 : tab2 = 23'b01110011110111100100000;
12'd1976 : tab2 = 23'b01110011101110101100000;
12'd1977 : tab2 = 23'b01110011100101110100111;
12'd1978 : tab2 = 23'b01110011011100111101101;
12'd1979 : tab2 = 23'b01110011010100000111010;
12'd1980 : tab2 = 23'b01110011001011010000111;
12'd1981 : tab2 = 23'b01110011000010011010101;
12'd1982 : tab2 = 23'b01110010111001100101001;
12'd1983 : tab2 = 23'b01110010110000101111111;
12'd1984 : tab2 = 23'b01110010100111111011001;
12'd1985 : tab2 = 23'b01110010011111000110100;
12'd1986 : tab2 = 23'b01110010010110010010010;
12'd1987 : tab2 = 23'b01110010001101011111000;
12'd1988 : tab2 = 23'b01110010000100101011011;
12'd1989 : tab2 = 23'b01110001111011111000101;
12'd1990 : tab2 = 23'b01110001110011000101101;
12'd1991 : tab2 = 23'b01110001101010010010110;
12'd1992 : tab2 = 23'b01110001100001100000110;
12'd1993 : tab2 = 23'b01110001011000101111000;
12'd1994 : tab2 = 23'b01110001001111111101110;
12'd1995 : tab2 = 23'b01110001000111001100101;
12'd1996 : tab2 = 23'b01110000111110011100000;
12'd1997 : tab2 = 23'b01110000110101101011101;
12'd1998 : tab2 = 23'b01110000101100111011111;
12'd1999 : tab2 = 23'b01110000100100001100010;
12'd2000 : tab2 = 23'b01110000011011011100111;
12'd2001 : tab2 = 23'b01110000010010101101101;
12'd2002 : tab2 = 23'b01110000001001111111000;
12'd2003 : tab2 = 23'b01110000000001010000111;
12'd2004 : tab2 = 23'b01101111111000100010111;
12'd2005 : tab2 = 23'b01101111101111110101100;
12'd2006 : tab2 = 23'b01101111100111001000001;
12'd2007 : tab2 = 23'b01101111011110011011010;
12'd2008 : tab2 = 23'b01101111010101101110100;
12'd2009 : tab2 = 23'b01101111001101000010110;
12'd2010 : tab2 = 23'b01101111000100010110110;
12'd2011 : tab2 = 23'b01101110111011101011101;
12'd2012 : tab2 = 23'b01101110110011000000010;
12'd2013 : tab2 = 23'b01101110101010010101000;
12'd2014 : tab2 = 23'b01101110100001101010101;
12'd2015 : tab2 = 23'b01101110011001000000011;
12'd2016 : tab2 = 23'b01101110010000010111001;
12'd2017 : tab2 = 23'b01101110000111101101100;
12'd2018 : tab2 = 23'b01101101111111000100000;
12'd2019 : tab2 = 23'b01101101110110011011010;
12'd2020 : tab2 = 23'b01101101101101110011001;
12'd2021 : tab2 = 23'b01101101100101001010111;
12'd2022 : tab2 = 23'b01101101011100100011001;
12'd2023 : tab2 = 23'b01101101010011111011111;
12'd2024 : tab2 = 23'b01101101001011010100100;
12'd2025 : tab2 = 23'b01101101000010101101100;
12'd2026 : tab2 = 23'b01101100111010000111011;
12'd2027 : tab2 = 23'b01101100110001100001001;
12'd2028 : tab2 = 23'b01101100101000111011101;
12'd2029 : tab2 = 23'b01101100100000010110010;
12'd2030 : tab2 = 23'b01101100010111110001010;
12'd2031 : tab2 = 23'b01101100001111001100000;
12'd2032 : tab2 = 23'b01101100000110100111111;
12'd2033 : tab2 = 23'b01101011111110000011111;
12'd2034 : tab2 = 23'b01101011110101100000001;
12'd2035 : tab2 = 23'b01101011101100111100110;
12'd2036 : tab2 = 23'b01101011100100011001100;
12'd2037 : tab2 = 23'b01101011011011110110110;
12'd2038 : tab2 = 23'b01101011010011010100101;
12'd2039 : tab2 = 23'b01101011001010110010101;
12'd2040 : tab2 = 23'b01101011000010010000111;
12'd2041 : tab2 = 23'b01101010111001101111100;
12'd2042 : tab2 = 23'b01101010110001001110010;
12'd2043 : tab2 = 23'b01101010101000101101110;
12'd2044 : tab2 = 23'b01101010100000001101001;
12'd2045 : tab2 = 23'b01101010010111101101011;
12'd2046 : tab2 = 23'b01101010001111001101011;
12'd2047 : tab2 = 23'b01101010000110101110010;
12'd2048 : tab2 = 23'b01101001111001111111110;
12'd2049 : tab2 = 23'b01101001101001000011000;
12'd2050 : tab2 = 23'b01101001011000000111101;
12'd2051 : tab2 = 23'b01101001000111001101011;
12'd2052 : tab2 = 23'b01101000110110010100100;
12'd2053 : tab2 = 23'b01101000100101011100111;
12'd2054 : tab2 = 23'b01101000010100100111000;
12'd2055 : tab2 = 23'b01101000000011110001111;
12'd2056 : tab2 = 23'b01100111110010111110001;
12'd2057 : tab2 = 23'b01100111100010001011111;
12'd2058 : tab2 = 23'b01100111010001011011011;
12'd2059 : tab2 = 23'b01100111000000101011011;
12'd2060 : tab2 = 23'b01100110101111111101000;
12'd2061 : tab2 = 23'b01100110011111010000000;
12'd2062 : tab2 = 23'b01100110001110100100010;
12'd2063 : tab2 = 23'b01100101111101111001101;
12'd2064 : tab2 = 23'b01100101101101010000101;
12'd2065 : tab2 = 23'b01100101011100101000101;
12'd2066 : tab2 = 23'b01100101001100000001111;
12'd2067 : tab2 = 23'b01100100111011011100110;
12'd2068 : tab2 = 23'b01100100101010111000110;
12'd2069 : tab2 = 23'b01100100011010010101110;
12'd2070 : tab2 = 23'b01100100001001110100000;
12'd2071 : tab2 = 23'b01100011111001010100010;
12'd2072 : tab2 = 23'b01100011101000110101000;
12'd2073 : tab2 = 23'b01100011011000010111011;
12'd2074 : tab2 = 23'b01100011000111111010111;
12'd2075 : tab2 = 23'b01100010110111011111111;
12'd2076 : tab2 = 23'b01100010100111000101111;
12'd2077 : tab2 = 23'b01100010010110101101101;
12'd2078 : tab2 = 23'b01100010000110010110010;
12'd2079 : tab2 = 23'b01100001110110000000001;
12'd2080 : tab2 = 23'b01100001100101101011001;
12'd2081 : tab2 = 23'b01100001010101010111111;
12'd2082 : tab2 = 23'b01100001000101000101011;
12'd2083 : tab2 = 23'b01100000110100110100001;
12'd2084 : tab2 = 23'b01100000100100100100101;
12'd2085 : tab2 = 23'b01100000010100010110001;
12'd2086 : tab2 = 23'b01100000000100001000110;
12'd2087 : tab2 = 23'b01011111110011111100100;
12'd2088 : tab2 = 23'b01011111100011110001110;
12'd2089 : tab2 = 23'b01011111010011101000011;
12'd2090 : tab2 = 23'b01011111000011011111110;
12'd2091 : tab2 = 23'b01011110110011011000100;
12'd2092 : tab2 = 23'b01011110100011010010101;
12'd2093 : tab2 = 23'b01011110010011001110001;
12'd2094 : tab2 = 23'b01011110000011001010100;
12'd2095 : tab2 = 23'b01011101110011001000001;
12'd2096 : tab2 = 23'b01011101100011000111010;
12'd2097 : tab2 = 23'b01011101010011000111100;
12'd2098 : tab2 = 23'b01011101000011001001001;
12'd2099 : tab2 = 23'b01011100110011001011101;
12'd2100 : tab2 = 23'b01011100100011001111101;
12'd2101 : tab2 = 23'b01011100010011010100100;
12'd2102 : tab2 = 23'b01011100000011011010111;
12'd2103 : tab2 = 23'b01011011110011100010101;
12'd2104 : tab2 = 23'b01011011100011101011001;
12'd2105 : tab2 = 23'b01011011010011110100110;
12'd2106 : tab2 = 23'b01011011000100000000100;
12'd2107 : tab2 = 23'b01011010110100001100110;
12'd2108 : tab2 = 23'b01011010100100011010000;
12'd2109 : tab2 = 23'b01011010010100101000101;
12'd2110 : tab2 = 23'b01011010000100111000110;
12'd2111 : tab2 = 23'b01011001110101001010000;
12'd2112 : tab2 = 23'b01011001100101011100010;
12'd2113 : tab2 = 23'b01011001010101101111101;
12'd2114 : tab2 = 23'b01011001000110000100001;
12'd2115 : tab2 = 23'b01011000110110011010011;
12'd2116 : tab2 = 23'b01011000100110110001011;
12'd2117 : tab2 = 23'b01011000010111001001001;
12'd2118 : tab2 = 23'b01011000000111100010111;
12'd2119 : tab2 = 23'b01010111110111111101100;
12'd2120 : tab2 = 23'b01010111101000011001010;
12'd2121 : tab2 = 23'b01010111011000110101111;
12'd2122 : tab2 = 23'b01010111001001010100000;
12'd2123 : tab2 = 23'b01010110111001110011011;
12'd2124 : tab2 = 23'b01010110101010010011111;
12'd2125 : tab2 = 23'b01010110011010110101101;
12'd2126 : tab2 = 23'b01010110001011011000101;
12'd2127 : tab2 = 23'b01010101111011111100000;
12'd2128 : tab2 = 23'b01010101101100100001010;
12'd2129 : tab2 = 23'b01010101011101000111110;
12'd2130 : tab2 = 23'b01010101001101101111001;
12'd2131 : tab2 = 23'b01010100111110010111100;
12'd2132 : tab2 = 23'b01010100101111000001101;
12'd2133 : tab2 = 23'b01010100011111101100001;
12'd2134 : tab2 = 23'b01010100010000011000011;
12'd2135 : tab2 = 23'b01010100000001000101101;
12'd2136 : tab2 = 23'b01010011110001110100000;
12'd2137 : tab2 = 23'b01010011100010100011001;
12'd2138 : tab2 = 23'b01010011010011010011101;
12'd2139 : tab2 = 23'b01010011000100000101100;
12'd2140 : tab2 = 23'b01010010110100111000101;
12'd2141 : tab2 = 23'b01010010100101101100011;
12'd2142 : tab2 = 23'b01010010010110100001100;
12'd2143 : tab2 = 23'b01010010000111010111110;
12'd2144 : tab2 = 23'b01010001111000001111100;
12'd2145 : tab2 = 23'b01010001101001000111110;
12'd2146 : tab2 = 23'b01010001011010000001100;
12'd2147 : tab2 = 23'b01010001001010111100011;
12'd2148 : tab2 = 23'b01010000111011111000100;
12'd2149 : tab2 = 23'b01010000101100110101011;
12'd2150 : tab2 = 23'b01010000011101110011011;
12'd2151 : tab2 = 23'b01010000001110110011000;
12'd2152 : tab2 = 23'b01001111111111110011010;
12'd2153 : tab2 = 23'b01001111110000110100110;
12'd2154 : tab2 = 23'b01001111100001110111001;
12'd2155 : tab2 = 23'b01001111010010111011011;
12'd2156 : tab2 = 23'b01001111000011111111111;
12'd2157 : tab2 = 23'b01001110110101000101110;
12'd2158 : tab2 = 23'b01001110100110001100101;
12'd2159 : tab2 = 23'b01001110010111010100110;
12'd2160 : tab2 = 23'b01001110001000011110011;
12'd2161 : tab2 = 23'b01001101111001101000011;
12'd2162 : tab2 = 23'b01001101101010110011111;
12'd2163 : tab2 = 23'b01001101011100000000101;
12'd2164 : tab2 = 23'b01001101001101001110001;
12'd2165 : tab2 = 23'b01001100111110011100110;
12'd2166 : tab2 = 23'b01001100101111101100111;
12'd2167 : tab2 = 23'b01001100100000111101011;
12'd2168 : tab2 = 23'b01001100010010001111111;
12'd2169 : tab2 = 23'b01001100000011100010110;
12'd2170 : tab2 = 23'b01001011110100110110110;
12'd2171 : tab2 = 23'b01001011100110001100001;
12'd2172 : tab2 = 23'b01001011010111100010100;
12'd2173 : tab2 = 23'b01001011001000111001100;
12'd2174 : tab2 = 23'b01001010111010010010001;
12'd2175 : tab2 = 23'b01001010101011101011110;
12'd2176 : tab2 = 23'b01001010011101000110101;
12'd2177 : tab2 = 23'b01001010001110100010100;
12'd2178 : tab2 = 23'b01001001111111111111000;
12'd2179 : tab2 = 23'b01001001110001011100110;
12'd2180 : tab2 = 23'b01001001100010111011110;
12'd2181 : tab2 = 23'b01001001010100011011101;
12'd2182 : tab2 = 23'b01001001000101111100100;
12'd2183 : tab2 = 23'b01001000110111011110100;
12'd2184 : tab2 = 23'b01001000101001000010000;
12'd2185 : tab2 = 23'b01001000011010100110000;
12'd2186 : tab2 = 23'b01001000001100001011011;
12'd2187 : tab2 = 23'b01000111111101110010000;
12'd2188 : tab2 = 23'b01000111101111011000111;
12'd2189 : tab2 = 23'b01000111100001000001110;
12'd2190 : tab2 = 23'b01000111010010101010111;
12'd2191 : tab2 = 23'b01000111000100010101010;
12'd2192 : tab2 = 23'b01000110110110000001011;
12'd2193 : tab2 = 23'b01000110100111101101101;
12'd2194 : tab2 = 23'b01000110011001011011101;
12'd2195 : tab2 = 23'b01000110001011001010011;
12'd2196 : tab2 = 23'b01000101111100111001101;
12'd2197 : tab2 = 23'b01000101101110101010101;
12'd2198 : tab2 = 23'b01000101100000011100100;
12'd2199 : tab2 = 23'b01000101010010001111010;
12'd2200 : tab2 = 23'b01000101000100000011000;
12'd2201 : tab2 = 23'b01000100110101110111110;
12'd2202 : tab2 = 23'b01000100100111101110000;
12'd2203 : tab2 = 23'b01000100011001100100110;
12'd2204 : tab2 = 23'b01000100001011011100110;
12'd2205 : tab2 = 23'b01000011111101010110000;
12'd2206 : tab2 = 23'b01000011101111010000000;
12'd2207 : tab2 = 23'b01000011100001001011000;
12'd2208 : tab2 = 23'b01000011010011000111001;
12'd2209 : tab2 = 23'b01000011000101000100001;
12'd2210 : tab2 = 23'b01000010110111000010100;
12'd2211 : tab2 = 23'b01000010101001000001101;
12'd2212 : tab2 = 23'b01000010011011000001110;
12'd2213 : tab2 = 23'b01000010001101000010111;
12'd2214 : tab2 = 23'b01000001111111000100111;
12'd2215 : tab2 = 23'b01000001110001001000011;
12'd2216 : tab2 = 23'b01000001100011001100011;
12'd2217 : tab2 = 23'b01000001010101010001011;
12'd2218 : tab2 = 23'b01000001000111010111111;
12'd2219 : tab2 = 23'b01000000111001011110110;
12'd2220 : tab2 = 23'b01000000101011100111000;
12'd2221 : tab2 = 23'b01000000011101110000011;
12'd2222 : tab2 = 23'b01000000001111111010001;
12'd2223 : tab2 = 23'b01000000000010000101110;
12'd2224 : tab2 = 23'b00111111110100010001110;
12'd2225 : tab2 = 23'b00111111100110011110111;
12'd2226 : tab2 = 23'b00111111011000101101010;
12'd2227 : tab2 = 23'b00111111001010111100010;
12'd2228 : tab2 = 23'b00111110111101001100100;
12'd2229 : tab2 = 23'b00111110101111011101010;
12'd2230 : tab2 = 23'b00111110100001101111101;
12'd2231 : tab2 = 23'b00111110010100000010100;
12'd2232 : tab2 = 23'b00111110000110010110111;
12'd2233 : tab2 = 23'b00111101111000101011111;
12'd2234 : tab2 = 23'b00111101101011000001101;
12'd2235 : tab2 = 23'b00111101011101011000111;
12'd2236 : tab2 = 23'b00111101001111110001001;
12'd2237 : tab2 = 23'b00111101000010001001110;
12'd2238 : tab2 = 23'b00111100110100100011101;
12'd2239 : tab2 = 23'b00111100100110111110110;
12'd2240 : tab2 = 23'b00111100011001011010101;
12'd2241 : tab2 = 23'b00111100001011110111100;
12'd2242 : tab2 = 23'b00111011111110010101010;
12'd2243 : tab2 = 23'b00111011110000110100000;
12'd2244 : tab2 = 23'b00111011100011010011111;
12'd2245 : tab2 = 23'b00111011010101110100011;
12'd2246 : tab2 = 23'b00111011001000010110000;
12'd2247 : tab2 = 23'b00111010111010111000101;
12'd2248 : tab2 = 23'b00111010101101011100011;
12'd2249 : tab2 = 23'b00111010100000000001000;
12'd2250 : tab2 = 23'b00111010010010100110100;
12'd2251 : tab2 = 23'b00111010000101001100110;
12'd2252 : tab2 = 23'b00111001110111110100001;
12'd2253 : tab2 = 23'b00111001101010011100100;
12'd2254 : tab2 = 23'b00111001011101000110000;
12'd2255 : tab2 = 23'b00111001001111110000100;
12'd2256 : tab2 = 23'b00111001000010011011010;
12'd2257 : tab2 = 23'b00111000110101000111101;
12'd2258 : tab2 = 23'b00111000100111110100101;
12'd2259 : tab2 = 23'b00111000011010100010011;
12'd2260 : tab2 = 23'b00111000001101010001100;
12'd2261 : tab2 = 23'b00111000000000000001011;
12'd2262 : tab2 = 23'b00110111110010110010010;
12'd2263 : tab2 = 23'b00110111100101100100001;
12'd2264 : tab2 = 23'b00110111011000010110100;
12'd2265 : tab2 = 23'b00110111001011001010010;
12'd2266 : tab2 = 23'b00110110111101111111000;
12'd2267 : tab2 = 23'b00110110110000110100011;
12'd2268 : tab2 = 23'b00110110100011101011000;
12'd2269 : tab2 = 23'b00110110010110100010001;
12'd2270 : tab2 = 23'b00110110001001011010100;
12'd2271 : tab2 = 23'b00110101111100010011110;
12'd2272 : tab2 = 23'b00110101101111001101111;
12'd2273 : tab2 = 23'b00110101100010001000111;
12'd2274 : tab2 = 23'b00110101010101000100101;
12'd2275 : tab2 = 23'b00110101001000000001100;
12'd2276 : tab2 = 23'b00110100111010111111011;
12'd2277 : tab2 = 23'b00110100101101111110010;
12'd2278 : tab2 = 23'b00110100100000111110001;
12'd2279 : tab2 = 23'b00110100010011111110100;
12'd2280 : tab2 = 23'b00110100000110111111110;
12'd2281 : tab2 = 23'b00110011111010000010010;
12'd2282 : tab2 = 23'b00110011101101000101101;
12'd2283 : tab2 = 23'b00110011100000001001011;
12'd2284 : tab2 = 23'b00110011010011001110111;
12'd2285 : tab2 = 23'b00110011000110010100110;
12'd2286 : tab2 = 23'b00110010111001011011101;
12'd2287 : tab2 = 23'b00110010101100100011010;
12'd2288 : tab2 = 23'b00110010011111101011111;
12'd2289 : tab2 = 23'b00110010010010110101100;
12'd2290 : tab2 = 23'b00110010000110000000001;
12'd2291 : tab2 = 23'b00110001111001001011100;
12'd2292 : tab2 = 23'b00110001101100011000000;
12'd2293 : tab2 = 23'b00110001011111100100101;
12'd2294 : tab2 = 23'b00110001010010110011001;
12'd2295 : tab2 = 23'b00110001000110000001111;
12'd2296 : tab2 = 23'b00110000111001010001110;
12'd2297 : tab2 = 23'b00110000101100100010101;
12'd2298 : tab2 = 23'b00110000011111110100001;
12'd2299 : tab2 = 23'b00110000010011000110110;
12'd2300 : tab2 = 23'b00110000000110011010000;
12'd2301 : tab2 = 23'b00101111111001101110010;
12'd2302 : tab2 = 23'b00101111101101000011101;
12'd2303 : tab2 = 23'b00101111100000011001111;
12'd2304 : tab2 = 23'b00101111010011110000100;
12'd2305 : tab2 = 23'b00101111000111001000010;
12'd2306 : tab2 = 23'b00101110111010100000111;
12'd2307 : tab2 = 23'b00101110101101111010110;
12'd2308 : tab2 = 23'b00101110100001010100110;
12'd2309 : tab2 = 23'b00101110010100110000001;
12'd2310 : tab2 = 23'b00101110001000001100101;
12'd2311 : tab2 = 23'b00101101111011101001010;
12'd2312 : tab2 = 23'b00101101101111000111001;
12'd2313 : tab2 = 23'b00101101100010100110010;
12'd2314 : tab2 = 23'b00101101010110000101110;
12'd2315 : tab2 = 23'b00101101001001100110010;
12'd2316 : tab2 = 23'b00101100111101000111110;
12'd2317 : tab2 = 23'b00101100110000101001101;
12'd2318 : tab2 = 23'b00101100100100001101000;
12'd2319 : tab2 = 23'b00101100010111110000111;
12'd2320 : tab2 = 23'b00101100001011010101110;
12'd2321 : tab2 = 23'b00101011111110111010111;
12'd2322 : tab2 = 23'b00101011110010100001111;
12'd2323 : tab2 = 23'b00101011100110001001000;
12'd2324 : tab2 = 23'b00101011011001110001010;
12'd2325 : tab2 = 23'b00101011001101011010011;
12'd2326 : tab2 = 23'b00101011000001000100000;
12'd2327 : tab2 = 23'b00101010110100101111010;
12'd2328 : tab2 = 23'b00101010101000011010110;
12'd2329 : tab2 = 23'b00101010011100000111010;
12'd2330 : tab2 = 23'b00101010001111110100001;
12'd2331 : tab2 = 23'b00101010000011100010011;
12'd2332 : tab2 = 23'b00101001110111010001010;
12'd2333 : tab2 = 23'b00101001101011000001001;
12'd2334 : tab2 = 23'b00101001011110110001101;
12'd2335 : tab2 = 23'b00101001010010100011100;
12'd2336 : tab2 = 23'b00101001000110010101110;
12'd2337 : tab2 = 23'b00101000111010001000111;
12'd2338 : tab2 = 23'b00101000101101111101000;
12'd2339 : tab2 = 23'b00101000100001110001101;
12'd2340 : tab2 = 23'b00101000010101100111011;
12'd2341 : tab2 = 23'b00101000001001011110010;
12'd2342 : tab2 = 23'b00100111111101010101011;
12'd2343 : tab2 = 23'b00100111110001001101100;
12'd2344 : tab2 = 23'b00100111100101000110010;
12'd2345 : tab2 = 23'b00100111011001000000011;
12'd2346 : tab2 = 23'b00100111001100111010111;
12'd2347 : tab2 = 23'b00100111000000110110100;
12'd2348 : tab2 = 23'b00100110110100110010101;
12'd2349 : tab2 = 23'b00100110101000101111110;
12'd2350 : tab2 = 23'b00100110011100101101110;
12'd2351 : tab2 = 23'b00100110010000101100011;
12'd2352 : tab2 = 23'b00100110000100101100001;
12'd2353 : tab2 = 23'b00100101111000101100011;
12'd2354 : tab2 = 23'b00100101101100101101110;
12'd2355 : tab2 = 23'b00100101100000101111011;
12'd2356 : tab2 = 23'b00100101010100110010101;
12'd2357 : tab2 = 23'b00100101001000110110001;
12'd2358 : tab2 = 23'b00100100111100111010110;
12'd2359 : tab2 = 23'b00100100110000111111101;
12'd2360 : tab2 = 23'b00100100100101000101111;
12'd2361 : tab2 = 23'b00100100011001001100011;
12'd2362 : tab2 = 23'b00100100001101010100001;
12'd2363 : tab2 = 23'b00100100000001011100111;
12'd2364 : tab2 = 23'b00100011110101100110000;
12'd2365 : tab2 = 23'b00100011101001110000000;
12'd2366 : tab2 = 23'b00100011011101111011001;
12'd2367 : tab2 = 23'b00100011010010000110011;
12'd2368 : tab2 = 23'b00100011000110010011001;
12'd2369 : tab2 = 23'b00100010111010100000011;
12'd2370 : tab2 = 23'b00100010101110101110101;
12'd2371 : tab2 = 23'b00100010100010111101101;
12'd2372 : tab2 = 23'b00100010010111001101001;
12'd2373 : tab2 = 23'b00100010001011011101101;
12'd2374 : tab2 = 23'b00100001111111101110110;
12'd2375 : tab2 = 23'b00100001110100000000111;
12'd2376 : tab2 = 23'b00100001101000010011101;
12'd2377 : tab2 = 23'b00100001011100100111011;
12'd2378 : tab2 = 23'b00100001010000111011101;
12'd2379 : tab2 = 23'b00100001000101010001000;
12'd2380 : tab2 = 23'b00100000111001100110111;
12'd2381 : tab2 = 23'b00100000101101111101100;
12'd2382 : tab2 = 23'b00100000100010010101000;
12'd2383 : tab2 = 23'b00100000010110101101001;
12'd2384 : tab2 = 23'b00100000001011000110010;
12'd2385 : tab2 = 23'b00011111111111100000011;
12'd2386 : tab2 = 23'b00011111110011111010110;
12'd2387 : tab2 = 23'b00011111101000010110001;
12'd2388 : tab2 = 23'b00011111011100110010011;
12'd2389 : tab2 = 23'b00011111010001001111101;
12'd2390 : tab2 = 23'b00011111000101101101010;
12'd2391 : tab2 = 23'b00011110111010001011110;
12'd2392 : tab2 = 23'b00011110101110101011010;
12'd2393 : tab2 = 23'b00011110100011001011000;
12'd2394 : tab2 = 23'b00011110010111101011110;
12'd2395 : tab2 = 23'b00011110001100001101100;
12'd2396 : tab2 = 23'b00011110000000110000001;
12'd2397 : tab2 = 23'b00011101110101010011000;
12'd2398 : tab2 = 23'b00011101101001110110111;
12'd2399 : tab2 = 23'b00011101011110011011101;
12'd2400 : tab2 = 23'b00011101010011000000110;
12'd2401 : tab2 = 23'b00011101000111100111001;
12'd2402 : tab2 = 23'b00011100111100001101111;
12'd2403 : tab2 = 23'b00011100110000110101110;
12'd2404 : tab2 = 23'b00011100100101011110000;
12'd2405 : tab2 = 23'b00011100011010000111010;
12'd2406 : tab2 = 23'b00011100001110110001011;
12'd2407 : tab2 = 23'b00011100000011011100001;
12'd2408 : tab2 = 23'b00011011111000000111100;
12'd2409 : tab2 = 23'b00011011101100110011111;
12'd2410 : tab2 = 23'b00011011100001100000110;
12'd2411 : tab2 = 23'b00011011010110001110010;
12'd2412 : tab2 = 23'b00011011001010111100110;
12'd2413 : tab2 = 23'b00011010111111101100001;
12'd2414 : tab2 = 23'b00011010110100011100010;
12'd2415 : tab2 = 23'b00011010101001001100100;
12'd2416 : tab2 = 23'b00011010011101111110001;
12'd2417 : tab2 = 23'b00011010010010110000011;
12'd2418 : tab2 = 23'b00011010000111100011100;
12'd2419 : tab2 = 23'b00011001111100010111010;
12'd2420 : tab2 = 23'b00011001110001001011010;
12'd2421 : tab2 = 23'b00011001100110000000101;
12'd2422 : tab2 = 23'b00011001011010110110100;
12'd2423 : tab2 = 23'b00011001001111101101000;
12'd2424 : tab2 = 23'b00011001000100100100011;
12'd2425 : tab2 = 23'b00011000111001011100010;
12'd2426 : tab2 = 23'b00011000101110010101010;
12'd2427 : tab2 = 23'b00011000100011001111001;
12'd2428 : tab2 = 23'b00011000011000001001010;
12'd2429 : tab2 = 23'b00011000001101000100100;
12'd2430 : tab2 = 23'b00011000000010000000010;
12'd2431 : tab2 = 23'b00010111110110111100010;
12'd2432 : tab2 = 23'b00010111101011111001100;
12'd2433 : tab2 = 23'b00010111100000110111101;
12'd2434 : tab2 = 23'b00010111010101110110001;
12'd2435 : tab2 = 23'b00010111001010110101111;
12'd2436 : tab2 = 23'b00010110111111110101111;
12'd2437 : tab2 = 23'b00010110110100110110100;
12'd2438 : tab2 = 23'b00010110101001111000000;
12'd2439 : tab2 = 23'b00010110011110111010011;
12'd2440 : tab2 = 23'b00010110010011111101011;
12'd2441 : tab2 = 23'b00010110001001000001000;
12'd2442 : tab2 = 23'b00010101111110000101101;
12'd2443 : tab2 = 23'b00010101110011001010111;
12'd2444 : tab2 = 23'b00010101101000010000101;
12'd2445 : tab2 = 23'b00010101011101010111010;
12'd2446 : tab2 = 23'b00010101010010011110001;
12'd2447 : tab2 = 23'b00010101000111100110011;
12'd2448 : tab2 = 23'b00010100111100101110111;
12'd2449 : tab2 = 23'b00010100110001111000101;
12'd2450 : tab2 = 23'b00010100100111000010100;
12'd2451 : tab2 = 23'b00010100011100001101011;
12'd2452 : tab2 = 23'b00010100010001011000111;
12'd2453 : tab2 = 23'b00010100000110100101010;
12'd2454 : tab2 = 23'b00010011111011110010010;
12'd2455 : tab2 = 23'b00010011110000111111101;
12'd2456 : tab2 = 23'b00010011100110001110000;
12'd2457 : tab2 = 23'b00010011011011011101001;
12'd2458 : tab2 = 23'b00010011010000101100110;
12'd2459 : tab2 = 23'b00010011000101111101011;
12'd2460 : tab2 = 23'b00010010111011001110100;
12'd2461 : tab2 = 23'b00010010110000100000011;
12'd2462 : tab2 = 23'b00010010100101110010101;
12'd2463 : tab2 = 23'b00010010011011000110010;
12'd2464 : tab2 = 23'b00010010010000011010000;
12'd2465 : tab2 = 23'b00010010000101101110110;
12'd2466 : tab2 = 23'b00010001111011000100001;
12'd2467 : tab2 = 23'b00010001110000011010001;
12'd2468 : tab2 = 23'b00010001100101110000100;
12'd2469 : tab2 = 23'b00010001011011001000000;
12'd2470 : tab2 = 23'b00010001010000100000010;
12'd2471 : tab2 = 23'b00010001000101111000111;
12'd2472 : tab2 = 23'b00010000111011010010010;
12'd2473 : tab2 = 23'b00010000110000101100011;
12'd2474 : tab2 = 23'b00010000100110000111011;
12'd2475 : tab2 = 23'b00010000011011100010111;
12'd2476 : tab2 = 23'b00010000010000111111000;
12'd2477 : tab2 = 23'b00010000000110011100000;
12'd2478 : tab2 = 23'b00001111111011111001101;
12'd2479 : tab2 = 23'b00001111110001010111100;
12'd2480 : tab2 = 23'b00001111100110110110100;
12'd2481 : tab2 = 23'b00001111011100010110010;
12'd2482 : tab2 = 23'b00001111010001110110100;
12'd2483 : tab2 = 23'b00001111000111010111010;
12'd2484 : tab2 = 23'b00001110111100111001000;
12'd2485 : tab2 = 23'b00001110110010011011010;
12'd2486 : tab2 = 23'b00001110100111111110011;
12'd2487 : tab2 = 23'b00001110011101100010001;
12'd2488 : tab2 = 23'b00001110010011000110001;
12'd2489 : tab2 = 23'b00001110001000101011001;
12'd2490 : tab2 = 23'b00001101111110010000111;
12'd2491 : tab2 = 23'b00001101110011110111010;
12'd2492 : tab2 = 23'b00001101101001011110001;
12'd2493 : tab2 = 23'b00001101011111000101101;
12'd2494 : tab2 = 23'b00001101010100101110000;
12'd2495 : tab2 = 23'b00001101001010010111011;
12'd2496 : tab2 = 23'b00001101000000000000111;
12'd2497 : tab2 = 23'b00001100110101101011010;
12'd2498 : tab2 = 23'b00001100101011010110010;
12'd2499 : tab2 = 23'b00001100100001000001111;
12'd2500 : tab2 = 23'b00001100010110101110000;
12'd2501 : tab2 = 23'b00001100001100011011010;
12'd2502 : tab2 = 23'b00001100000010001000100;
12'd2503 : tab2 = 23'b00001011110111110110110;
12'd2504 : tab2 = 23'b00001011101101100101110;
12'd2505 : tab2 = 23'b00001011100011010101010;
12'd2506 : tab2 = 23'b00001011011001000101110;
12'd2507 : tab2 = 23'b00001011001110110110100;
12'd2508 : tab2 = 23'b00001011000100101000001;
12'd2509 : tab2 = 23'b00001010111010011010011;
12'd2510 : tab2 = 23'b00001010110000001101001;
12'd2511 : tab2 = 23'b00001010100110000000101;
12'd2512 : tab2 = 23'b00001010011011110100111;
12'd2513 : tab2 = 23'b00001010010001101001011;
12'd2514 : tab2 = 23'b00001010000111011110111;
12'd2515 : tab2 = 23'b00001001111101010100110;
12'd2516 : tab2 = 23'b00001001110011001011110;
12'd2517 : tab2 = 23'b00001001101001000011001;
12'd2518 : tab2 = 23'b00001001011110111011010;
12'd2519 : tab2 = 23'b00001001010100110011110;
12'd2520 : tab2 = 23'b00001001001010101101000;
12'd2521 : tab2 = 23'b00001001000000100110111;
12'd2522 : tab2 = 23'b00001000110110100001101;
12'd2523 : tab2 = 23'b00001000101100011100111;
12'd2524 : tab2 = 23'b00001000100010011000110;
12'd2525 : tab2 = 23'b00001000011000010101001;
12'd2526 : tab2 = 23'b00001000001110010010011;
12'd2527 : tab2 = 23'b00001000000100010000001;
12'd2528 : tab2 = 23'b00000111111010001110101;
12'd2529 : tab2 = 23'b00000111110000001101010;
12'd2530 : tab2 = 23'b00000111100110001101011;
12'd2531 : tab2 = 23'b00000111011100001101101;
12'd2532 : tab2 = 23'b00000111010010001110101;
12'd2533 : tab2 = 23'b00000111001000010000000;
12'd2534 : tab2 = 23'b00000110111110010010001;
12'd2535 : tab2 = 23'b00000110110100010101000;
12'd2536 : tab2 = 23'b00000110101010011000011;
12'd2537 : tab2 = 23'b00000110100000011100101;
12'd2538 : tab2 = 23'b00000110010110100001100;
12'd2539 : tab2 = 23'b00000110001100100110101;
12'd2540 : tab2 = 23'b00000110000010101100111;
12'd2541 : tab2 = 23'b00000101111000110011000;
12'd2542 : tab2 = 23'b00000101101110111010011;
12'd2543 : tab2 = 23'b00000101100101000010000;
12'd2544 : tab2 = 23'b00000101011011001010100;
12'd2545 : tab2 = 23'b00000101010001010011110;
12'd2546 : tab2 = 23'b00000101000111011101011;
12'd2547 : tab2 = 23'b00000100111101100111110;
12'd2548 : tab2 = 23'b00000100110011110010101;
12'd2549 : tab2 = 23'b00000100101001111110100;
12'd2550 : tab2 = 23'b00000100100000001010001;
12'd2551 : tab2 = 23'b00000100010110010111011;
12'd2552 : tab2 = 23'b00000100001100100100100;
12'd2553 : tab2 = 23'b00000100000010110010100;
12'd2554 : tab2 = 23'b00000011111001000001000;
12'd2555 : tab2 = 23'b00000011101111010000100;
12'd2556 : tab2 = 23'b00000011100101100000001;
12'd2557 : tab2 = 23'b00000011011011110000100;
12'd2558 : tab2 = 23'b00000011010010000001111;
12'd2559 : tab2 = 23'b00000011001000010011011;
12'd2560 : tab2 = 23'b00000010111110100101110;
12'd2561 : tab2 = 23'b00000010110100111000100;
12'd2562 : tab2 = 23'b00000010101011001100000;
12'd2563 : tab2 = 23'b00000010100001100000010;
12'd2564 : tab2 = 23'b00000010010111110100111;
12'd2565 : tab2 = 23'b00000010001110001010010;
12'd2566 : tab2 = 23'b00000010000100011111111;
12'd2567 : tab2 = 23'b00000001111010110110011;
12'd2568 : tab2 = 23'b00000001110001001101011;
12'd2569 : tab2 = 23'b00000001100111100101010;
12'd2570 : tab2 = 23'b00000001011101111101101;
12'd2571 : tab2 = 23'b00000001010100010110101;
12'd2572 : tab2 = 23'b00000001001010101111111;
12'd2573 : tab2 = 23'b00000001000001001010001;
12'd2574 : tab2 = 23'b00000000110111100100101;
12'd2575 : tab2 = 23'b00000000101110000000000;
12'd2576 : tab2 = 23'b00000000100100011100000;
12'd2577 : tab2 = 23'b00000000011010111000100;
12'd2578 : tab2 = 23'b00000000010001010101011;
12'd2579 : tab2 = 23'b00000000000111110011000;
12'd2580 : tab2 = 23'b11111111111100100010101;
12'd2581 : tab2 = 23'b11111111101001100000100;
12'd2582 : tab2 = 23'b11111111010110011111011;
12'd2583 : tab2 = 23'b11111111000011011111011;
12'd2584 : tab2 = 23'b11111110110000100000010;
12'd2585 : tab2 = 23'b11111110011101100010111;
12'd2586 : tab2 = 23'b11111110001010100110100;
12'd2587 : tab2 = 23'b11111101110111101010110;
12'd2588 : tab2 = 23'b11111101100100110001001;
12'd2589 : tab2 = 23'b11111101010001111000000;
12'd2590 : tab2 = 23'b11111100111111000000110;
12'd2591 : tab2 = 23'b11111100101100001001110;
12'd2592 : tab2 = 23'b11111100011001010100011;
12'd2593 : tab2 = 23'b11111100000110100000001;
12'd2594 : tab2 = 23'b11111011110011101100111;
12'd2595 : tab2 = 23'b11111011100000111010110;
12'd2596 : tab2 = 23'b11111011001110001010001;
12'd2597 : tab2 = 23'b11111010111011011010001;
12'd2598 : tab2 = 23'b11111010101000101100010;
12'd2599 : tab2 = 23'b11111010010101111110111;
12'd2600 : tab2 = 23'b11111010000011010010101;
12'd2601 : tab2 = 23'b11111001110000101000000;
12'd2602 : tab2 = 23'b11111001011101111101110;
12'd2603 : tab2 = 23'b11111001001011010101001;
12'd2604 : tab2 = 23'b11111000111000101101101;
12'd2605 : tab2 = 23'b11111000100110000111010;
12'd2606 : tab2 = 23'b11111000010011100001001;
12'd2607 : tab2 = 23'b11111000000000111101011;
12'd2608 : tab2 = 23'b11110111101110011010000;
12'd2609 : tab2 = 23'b11110111011011111000010;
12'd2610 : tab2 = 23'b11110111001001010111110;
12'd2611 : tab2 = 23'b11110110110110111000001;
12'd2612 : tab2 = 23'b11110110100100011001011;
12'd2613 : tab2 = 23'b11110110010001111011111;
12'd2614 : tab2 = 23'b11110101111111100000000;
12'd2615 : tab2 = 23'b11110101101101000100101;
12'd2616 : tab2 = 23'b11110101011010101010110;
12'd2617 : tab2 = 23'b11110101001000010010000;
12'd2618 : tab2 = 23'b11110100110101111010010;
12'd2619 : tab2 = 23'b11110100100011100011100;
12'd2620 : tab2 = 23'b11110100010001001101110;
12'd2621 : tab2 = 23'b11110011111110111001110;
12'd2622 : tab2 = 23'b11110011101100100110101;
12'd2623 : tab2 = 23'b11110011011010010100000;
12'd2624 : tab2 = 23'b11110011001000000011101;
12'd2625 : tab2 = 23'b11110010110101110011110;
12'd2626 : tab2 = 23'b11110010100011100100111;
12'd2627 : tab2 = 23'b11110010010001010111011;
12'd2628 : tab2 = 23'b11110001111111001010101;
12'd2629 : tab2 = 23'b11110001101100111111011;
12'd2630 : tab2 = 23'b11110001011010110100000;
12'd2631 : tab2 = 23'b11110001001000101011011;
12'd2632 : tab2 = 23'b11110000110110100011010;
12'd2633 : tab2 = 23'b11110000100100011100101;
12'd2634 : tab2 = 23'b11110000010010010110101;
12'd2635 : tab2 = 23'b11110000000000010000111;
12'd2636 : tab2 = 23'b11101111101110001101111;
12'd2637 : tab2 = 23'b11101111011100001011100;
12'd2638 : tab2 = 23'b11101111001010001001011;
12'd2639 : tab2 = 23'b11101110111000001001000;
12'd2640 : tab2 = 23'b11101110100110001001101;
12'd2641 : tab2 = 23'b11101110010100001011110;
12'd2642 : tab2 = 23'b11101110000010001101110;
12'd2643 : tab2 = 23'b11101101110000010010000;
12'd2644 : tab2 = 23'b11101101011110010110101;
12'd2645 : tab2 = 23'b11101101001100011101011;
12'd2646 : tab2 = 23'b11101100111010100011100;
12'd2647 : tab2 = 23'b11101100101000101100011;
12'd2648 : tab2 = 23'b11101100010110110101110;
12'd2649 : tab2 = 23'b11101100000101000000000;
12'd2650 : tab2 = 23'b11101011110011001011111;
12'd2651 : tab2 = 23'b11101011100001011000001;
12'd2652 : tab2 = 23'b11101011001111100101011;
12'd2653 : tab2 = 23'b11101010111101110011110;
12'd2654 : tab2 = 23'b11101010101100000100010;
12'd2655 : tab2 = 23'b11101010011010010101011;
12'd2656 : tab2 = 23'b11101010001000100110101;
12'd2657 : tab2 = 23'b11101001110110111001100;
12'd2658 : tab2 = 23'b11101001100101001101100;
12'd2659 : tab2 = 23'b11101001010011100011000;
12'd2660 : tab2 = 23'b11101001000001111000111;
12'd2661 : tab2 = 23'b11101000110000010000100;
12'd2662 : tab2 = 23'b11101000011110100111110;
12'd2663 : tab2 = 23'b11101000001101000001011;
12'd2664 : tab2 = 23'b11100111111011011011111;
12'd2665 : tab2 = 23'b11100111101001110111011;
12'd2666 : tab2 = 23'b11100111011000010100000;
12'd2667 : tab2 = 23'b11100111000110110001011;
12'd2668 : tab2 = 23'b11100110110101010000000;
12'd2669 : tab2 = 23'b11100110100011101111100;
12'd2670 : tab2 = 23'b11100110010010001111111;
12'd2671 : tab2 = 23'b11100110000000110010000;
12'd2672 : tab2 = 23'b11100101101111010100100;
12'd2673 : tab2 = 23'b11100101011101111000101;
12'd2674 : tab2 = 23'b11100101001100011101101;
12'd2675 : tab2 = 23'b11100100111011000011000;
12'd2676 : tab2 = 23'b11100100101001101010001;
12'd2677 : tab2 = 23'b11100100011000010010001;
12'd2678 : tab2 = 23'b11100100000110111011001;
12'd2679 : tab2 = 23'b11100011110101100101001;
12'd2680 : tab2 = 23'b11100011100100010000110;
12'd2681 : tab2 = 23'b11100011010010111100110;
12'd2682 : tab2 = 23'b11100011000001101010001;
12'd2683 : tab2 = 23'b11100010110000011000001;
12'd2684 : tab2 = 23'b11100010011111000111110;
12'd2685 : tab2 = 23'b11100010001101110111100;
12'd2686 : tab2 = 23'b11100001111100101001000;
12'd2687 : tab2 = 23'b11100001101011011011000;
12'd2688 : tab2 = 23'b11100001011010001110011;
12'd2689 : tab2 = 23'b11100001001001000010110;
12'd2690 : tab2 = 23'b11100000110111110111100;
12'd2691 : tab2 = 23'b11100000100110101110100;
12'd2692 : tab2 = 23'b11100000010101100101111;
12'd2693 : tab2 = 23'b11100000000100011110010;
12'd2694 : tab2 = 23'b11011111110011011000000;
12'd2695 : tab2 = 23'b11011111100010010001110;
12'd2696 : tab2 = 23'b11011111010001001110001;
12'd2697 : tab2 = 23'b11011111000000001010011;
12'd2698 : tab2 = 23'b11011110101111000111101;
12'd2699 : tab2 = 23'b11011110011110000101101;
12'd2700 : tab2 = 23'b11011110001101000110000;
12'd2701 : tab2 = 23'b11011101111100000110101;
12'd2702 : tab2 = 23'b11011101101011000111110;
12'd2703 : tab2 = 23'b11011101011010001010100;
12'd2704 : tab2 = 23'b11011101001001001101011;
12'd2705 : tab2 = 23'b11011100111000010010000;
12'd2706 : tab2 = 23'b11011100100111011000000;
12'd2707 : tab2 = 23'b11011100010110011110101;
12'd2708 : tab2 = 23'b11011100000101100101100;
12'd2709 : tab2 = 23'b11011011110100101110100;
12'd2710 : tab2 = 23'b11011011100011110111111;
12'd2711 : tab2 = 23'b11011011010011000010010;
12'd2712 : tab2 = 23'b11011011000010001110001;
12'd2713 : tab2 = 23'b11011010110001011010100;
12'd2714 : tab2 = 23'b11011010100000101000011;
12'd2715 : tab2 = 23'b11011010001111110110100;
12'd2716 : tab2 = 23'b11011001111111000110010;
12'd2717 : tab2 = 23'b11011001101110010110010;
12'd2718 : tab2 = 23'b11011001011101101000000;
12'd2719 : tab2 = 23'b11011001001100111010001;
12'd2720 : tab2 = 23'b11011000111100001101110;
12'd2721 : tab2 = 23'b11011000101011100010001;
12'd2722 : tab2 = 23'b11011000011010110111001;
12'd2723 : tab2 = 23'b11011000001010001110001;
12'd2724 : tab2 = 23'b11010111111001100101101;
12'd2725 : tab2 = 23'b11010111101000111101011;
12'd2726 : tab2 = 23'b11010111011000010110101;
12'd2727 : tab2 = 23'b11010111000111110001011;
12'd2728 : tab2 = 23'b11010110110111001100101;
12'd2729 : tab2 = 23'b11010110100110101000010;
12'd2730 : tab2 = 23'b11010110010110000101100;
12'd2731 : tab2 = 23'b11010110000101100100000;
12'd2732 : tab2 = 23'b11010101110101000011000;
12'd2733 : tab2 = 23'b11010101100100100011000;
12'd2734 : tab2 = 23'b11010101010100000100011;
12'd2735 : tab2 = 23'b11010101000011100110010;
12'd2736 : tab2 = 23'b11010100110011001001110;
12'd2737 : tab2 = 23'b11010100100010101100111;
12'd2738 : tab2 = 23'b11010100010010010001101;
12'd2739 : tab2 = 23'b11010100000001110111110;
12'd2740 : tab2 = 23'b11010011110001011110011;
12'd2741 : tab2 = 23'b11010011100001000110100;
12'd2742 : tab2 = 23'b11010011010000101111000;
12'd2743 : tab2 = 23'b11010011000000011001000;
12'd2744 : tab2 = 23'b11010010110000000011010;
12'd2745 : tab2 = 23'b11010010011111101111001;
12'd2746 : tab2 = 23'b11010010001111011011011;
12'd2747 : tab2 = 23'b11010001111111001001001;
12'd2748 : tab2 = 23'b11010001101110110111010;
12'd2749 : tab2 = 23'b11010001011110100110111;
12'd2750 : tab2 = 23'b11010001001110010110111;
12'd2751 : tab2 = 23'b11010000111110001000011;
12'd2752 : tab2 = 23'b11010000101101111010001;
12'd2753 : tab2 = 23'b11010000011101101101100;
12'd2754 : tab2 = 23'b11010000001101100001110;
12'd2755 : tab2 = 23'b11001111111101010110100;
12'd2756 : tab2 = 23'b11001111101101001100101;
12'd2757 : tab2 = 23'b11001111011101000011101;
12'd2758 : tab2 = 23'b11001111001100111011110;
12'd2759 : tab2 = 23'b11001110111100110100110;
12'd2760 : tab2 = 23'b11001110101100101110000;
12'd2761 : tab2 = 23'b11001110011100101000110;
12'd2762 : tab2 = 23'b11001110001100100100000;
12'd2763 : tab2 = 23'b11001101111100100000101;
12'd2764 : tab2 = 23'b11001101101100011110010;
12'd2765 : tab2 = 23'b11001101011100011100001;
12'd2766 : tab2 = 23'b11001101001100011100001;
12'd2767 : tab2 = 23'b11001100111100011100100;
12'd2768 : tab2 = 23'b11001100101100011101011;
12'd2769 : tab2 = 23'b11001100011100011111100;
12'd2770 : tab2 = 23'b11001100001100100010000;
12'd2771 : tab2 = 23'b11001011111100100110001;
12'd2772 : tab2 = 23'b11001011101100101010101;
12'd2773 : tab2 = 23'b11001011011100110000100;
12'd2774 : tab2 = 23'b11001011001100110111011;
12'd2775 : tab2 = 23'b11001010111100111110100;
12'd2776 : tab2 = 23'b11001010101101000111110;
12'd2777 : tab2 = 23'b11001010011101010000010;
12'd2778 : tab2 = 23'b11001010001101011011010;
12'd2779 : tab2 = 23'b11001001111101100110001;
12'd2780 : tab2 = 23'b11001001101101110010100;
12'd2781 : tab2 = 23'b11001001011101111111111;
12'd2782 : tab2 = 23'b11001001001110001101100;
12'd2783 : tab2 = 23'b11001000111110011100100;
12'd2784 : tab2 = 23'b11001000101110101100000;
12'd2785 : tab2 = 23'b11001000011110111100111;
12'd2786 : tab2 = 23'b11001000001111001110001;
12'd2787 : tab2 = 23'b11000111111111100000111;
12'd2788 : tab2 = 23'b11000111101111110011111;
12'd2789 : tab2 = 23'b11000111100000001000100;
12'd2790 : tab2 = 23'b11000111010000011101011;
12'd2791 : tab2 = 23'b11000111000000110011110;
12'd2792 : tab2 = 23'b11000110110001001010101;
12'd2793 : tab2 = 23'b11000110100001100010110;
12'd2794 : tab2 = 23'b11000110010001111011010;
12'd2795 : tab2 = 23'b11000110000010010101010;
12'd2796 : tab2 = 23'b11000101110010101111101;
12'd2797 : tab2 = 23'b11000101100011001011100;
12'd2798 : tab2 = 23'b11000101010011100111101;
12'd2799 : tab2 = 23'b11000101000100000100110;
12'd2800 : tab2 = 23'b11000100110100100010110;
12'd2801 : tab2 = 23'b11000100100101000010001;
12'd2802 : tab2 = 23'b11000100010101100001100;
12'd2803 : tab2 = 23'b11000100000110000010001;
12'd2804 : tab2 = 23'b11000011110110100100010;
12'd2805 : tab2 = 23'b11000011100111000110110;
12'd2806 : tab2 = 23'b11000011010111101010001;
12'd2807 : tab2 = 23'b11000011001000001110011;
12'd2808 : tab2 = 23'b11000010111000110011110;
12'd2809 : tab2 = 23'b11000010101001011001110;
12'd2810 : tab2 = 23'b11000010011010000000010;
12'd2811 : tab2 = 23'b11000010001010101000101;
12'd2812 : tab2 = 23'b11000001111011010001011;
12'd2813 : tab2 = 23'b11000001101011111010100;
12'd2814 : tab2 = 23'b11000001011100100101010;
12'd2815 : tab2 = 23'b11000001001101010000001;
12'd2816 : tab2 = 23'b11000000111101111100100;
12'd2817 : tab2 = 23'b11000000101110101001110;
12'd2818 : tab2 = 23'b11000000011111010111011;
12'd2819 : tab2 = 23'b11000000010000000110010;
12'd2820 : tab2 = 23'b11000000000000110101101;
12'd2821 : tab2 = 23'b10111111110001100110000;
12'd2822 : tab2 = 23'b10111111100010010111110;
12'd2823 : tab2 = 23'b10111111010011001001110;
12'd2824 : tab2 = 23'b10111111000011111101010;
12'd2825 : tab2 = 23'b10111110110100110001001;
12'd2826 : tab2 = 23'b10111110100101100101111;
12'd2827 : tab2 = 23'b10111110010110011100000;
12'd2828 : tab2 = 23'b10111110000111010001111;
12'd2829 : tab2 = 23'b10111101111000001001011;
12'd2830 : tab2 = 23'b10111101101001000010001;
12'd2831 : tab2 = 23'b10111101011001111010110;
12'd2832 : tab2 = 23'b10111101001010110100110;
12'd2833 : tab2 = 23'b10111100111011101111101;
12'd2834 : tab2 = 23'b10111100101100101010111;
12'd2835 : tab2 = 23'b10111100011101100111101;
12'd2836 : tab2 = 23'b10111100001110100101001;
12'd2837 : tab2 = 23'b10111011111111100011001;
12'd2838 : tab2 = 23'b10111011110000100010111;
12'd2839 : tab2 = 23'b10111011100001100010001;
12'd2840 : tab2 = 23'b10111011010010100010101;
12'd2841 : tab2 = 23'b10111011000011100100100;
12'd2842 : tab2 = 23'b10111010110100100110111;
12'd2843 : tab2 = 23'b10111010100101101010101;
12'd2844 : tab2 = 23'b10111010010110101110101;
12'd2845 : tab2 = 23'b10111010000111110011000;
12'd2846 : tab2 = 23'b10111001111000111000111;
12'd2847 : tab2 = 23'b10111001101010000000000;
12'd2848 : tab2 = 23'b10111001011011000111100;
12'd2849 : tab2 = 23'b10111001001100001111011;
12'd2850 : tab2 = 23'b10111000111101011000110;
12'd2851 : tab2 = 23'b10111000101110100010011;
12'd2852 : tab2 = 23'b10111000011111101101011;
12'd2853 : tab2 = 23'b10111000010000111000111;
12'd2854 : tab2 = 23'b10111000000010000101101;
12'd2855 : tab2 = 23'b10110111110011010010101;
12'd2856 : tab2 = 23'b10110111100100100001010;
12'd2857 : tab2 = 23'b10110111010101110000001;
12'd2858 : tab2 = 23'b10110111000110111111110;
12'd2859 : tab2 = 23'b10110110111000010000011;
12'd2860 : tab2 = 23'b10110110101001100001111;
12'd2861 : tab2 = 23'b10110110011010110100001;
12'd2862 : tab2 = 23'b10110110001100000110111;
12'd2863 : tab2 = 23'b10110101111101011010111;
12'd2864 : tab2 = 23'b10110101101110101111111;
12'd2865 : tab2 = 23'b10110101100000000101000;
12'd2866 : tab2 = 23'b10110101010001011011001;
12'd2867 : tab2 = 23'b10110101000010110010100;
12'd2868 : tab2 = 23'b10110100110100001010100;
12'd2869 : tab2 = 23'b10110100100101100011101;
12'd2870 : tab2 = 23'b10110100010110111101001;
12'd2871 : tab2 = 23'b10110100001000010111110;
12'd2872 : tab2 = 23'b10110011111001110010011;
12'd2873 : tab2 = 23'b10110011101011001111001;
12'd2874 : tab2 = 23'b10110011011100101100001;
12'd2875 : tab2 = 23'b10110011001110001001011;
12'd2876 : tab2 = 23'b10110010111111101000001;
12'd2877 : tab2 = 23'b10110010110001000111001;
12'd2878 : tab2 = 23'b10110010100010100111100;
12'd2879 : tab2 = 23'b10110010010100001000010;
12'd2880 : tab2 = 23'b10110010000101101001111;
12'd2881 : tab2 = 23'b10110001110111001100011;
12'd2882 : tab2 = 23'b10110001101000101111101;
12'd2883 : tab2 = 23'b10110001011010010011111;
12'd2884 : tab2 = 23'b10110001001011111000111;
12'd2885 : tab2 = 23'b10110000111101011110001;
12'd2886 : tab2 = 23'b10110000101111000100111;
12'd2887 : tab2 = 23'b10110000100000101011111;
12'd2888 : tab2 = 23'b10110000010010010011111;
12'd2889 : tab2 = 23'b10110000000011111101001;
12'd2890 : tab2 = 23'b10101111110101100110101;
12'd2891 : tab2 = 23'b10101111100111010001001;
12'd2892 : tab2 = 23'b10101111011000111100111;
12'd2893 : tab2 = 23'b10101111001010101000101;
12'd2894 : tab2 = 23'b10101110111100010101100;
12'd2895 : tab2 = 23'b10101110101110000010110;
12'd2896 : tab2 = 23'b10101110011111110001011;
12'd2897 : tab2 = 23'b10101110010001100001001;
12'd2898 : tab2 = 23'b10101110000011010000111;
12'd2899 : tab2 = 23'b10101101110101000001101;
12'd2900 : tab2 = 23'b10101101100110110011101;
12'd2901 : tab2 = 23'b10101101011000100101111;
12'd2902 : tab2 = 23'b10101101001010011000101;
12'd2903 : tab2 = 23'b10101100111100001100101;
12'd2904 : tab2 = 23'b10101100101110000001101;
12'd2905 : tab2 = 23'b10101100011111110110110;
12'd2906 : tab2 = 23'b10101100010001101101011;
12'd2907 : tab2 = 23'b10101100000011100100010;
12'd2908 : tab2 = 23'b10101011110101011011111;
12'd2909 : tab2 = 23'b10101011100111010101000;
12'd2910 : tab2 = 23'b10101011011001001110011;
12'd2911 : tab2 = 23'b10101011001011001000010;
12'd2912 : tab2 = 23'b10101010111101000011010;
12'd2913 : tab2 = 23'b10101010101110111111001;
12'd2914 : tab2 = 23'b10101010100000111011010;
12'd2915 : tab2 = 23'b10101010010010111000111;
12'd2916 : tab2 = 23'b10101010000100110110111;
12'd2917 : tab2 = 23'b10101001110110110101100;
12'd2918 : tab2 = 23'b10101001101000110101001;
12'd2919 : tab2 = 23'b10101001011010110101101;
12'd2920 : tab2 = 23'b10101001001100110110110;
12'd2921 : tab2 = 23'b10101000111110111000110;
12'd2922 : tab2 = 23'b10101000110000111011010;
12'd2923 : tab2 = 23'b10101000100010111111000;
12'd2924 : tab2 = 23'b10101000010101000010111;
12'd2925 : tab2 = 23'b10101000000111000111011;
12'd2926 : tab2 = 23'b10100111111001001100111;
12'd2927 : tab2 = 23'b10100111101011010011100;
12'd2928 : tab2 = 23'b10100111011101011010111;
12'd2929 : tab2 = 23'b10100111001111100011000;
12'd2930 : tab2 = 23'b10100111000001101011011;
12'd2931 : tab2 = 23'b10100110110011110101010;
12'd2932 : tab2 = 23'b10100110100101111111011;
12'd2933 : tab2 = 23'b10100110011000001010011;
12'd2934 : tab2 = 23'b10100110001010010110001;
12'd2935 : tab2 = 23'b10100101111100100010110;
12'd2936 : tab2 = 23'b10100101101110101111110;
12'd2937 : tab2 = 23'b10100101100000111110000;
12'd2938 : tab2 = 23'b10100101010011001100011;
12'd2939 : tab2 = 23'b10100101000101011100011;
12'd2940 : tab2 = 23'b10100100110111101100101;
12'd2941 : tab2 = 23'b10100100101001111101000;
12'd2942 : tab2 = 23'b10100100011100001110111;
12'd2943 : tab2 = 23'b10100100001110100001100;
12'd2944 : tab2 = 23'b10100100000000110100100;
12'd2945 : tab2 = 23'b10100011110011001000010;
12'd2946 : tab2 = 23'b10100011100101011101011;
12'd2947 : tab2 = 23'b10100011010111110010111;
12'd2948 : tab2 = 23'b10100011001010001001000;
12'd2949 : tab2 = 23'b10100010111100100000001;
12'd2950 : tab2 = 23'b10100010101110110111100;
12'd2951 : tab2 = 23'b10100010100001010000000;
12'd2952 : tab2 = 23'b10100010010011101001101;
12'd2953 : tab2 = 23'b10100010000110000010111;
12'd2954 : tab2 = 23'b10100001111000011101011;
12'd2955 : tab2 = 23'b10100001101010111001000;
12'd2956 : tab2 = 23'b10100001011101010101001;
12'd2957 : tab2 = 23'b10100001001111110010001;
12'd2958 : tab2 = 23'b10100001000010001111100;
12'd2959 : tab2 = 23'b10100000110100101110010;
12'd2960 : tab2 = 23'b10100000100111001100101;
12'd2961 : tab2 = 23'b10100000011001101100111;
12'd2962 : tab2 = 23'b10100000001100001101100;
12'd2963 : tab2 = 23'b10011111111110101110011;
12'd2964 : tab2 = 23'b10011111110001010000101;
12'd2965 : tab2 = 23'b10011111100011110011001;
12'd2966 : tab2 = 23'b10011111010110010110111;
12'd2967 : tab2 = 23'b10011111001000111010011;
12'd2968 : tab2 = 23'b10011110111011011111011;
12'd2969 : tab2 = 23'b10011110101110000101001;
12'd2970 : tab2 = 23'b10011110100000101011001;
12'd2971 : tab2 = 23'b10011110010011010010000;
12'd2972 : tab2 = 23'b10011110000101111010001;
12'd2973 : tab2 = 23'b10011101111000100010100;
12'd2974 : tab2 = 23'b10011101101011001011001;
12'd2975 : tab2 = 23'b10011101011101110101010;
12'd2976 : tab2 = 23'b10011101010000100000000;
12'd2977 : tab2 = 23'b10011101000011001011001;
12'd2978 : tab2 = 23'b10011100110101110111010;
12'd2979 : tab2 = 23'b10011100101000100100011;
12'd2980 : tab2 = 23'b10011100011011010001111;
12'd2981 : tab2 = 23'b10011100001101111111110;
12'd2982 : tab2 = 23'b10011100000000101110111;
12'd2983 : tab2 = 23'b10011011110011011110011;
12'd2984 : tab2 = 23'b10011011100110001111000;
12'd2985 : tab2 = 23'b10011011011001000000001;
12'd2986 : tab2 = 23'b10011011001011110001011;
12'd2987 : tab2 = 23'b10011010111110100100000;
12'd2988 : tab2 = 23'b10011010110001010110111;
12'd2989 : tab2 = 23'b10011010100100001011001;
12'd2990 : tab2 = 23'b10011010010110111111100;
12'd2991 : tab2 = 23'b10011010001001110100010;
12'd2992 : tab2 = 23'b10011001111100101010011;
12'd2993 : tab2 = 23'b10011001101111100001110;
12'd2994 : tab2 = 23'b10011001100010011000011;
12'd2995 : tab2 = 23'b10011001010101010000111;
12'd2996 : tab2 = 23'b10011001001000001001100;
12'd2997 : tab2 = 23'b10011000111011000011000;
12'd2998 : tab2 = 23'b10011000101101111101011;
12'd2999 : tab2 = 23'b10011000100000111000001;
12'd3000 : tab2 = 23'b10011000010011110011011;
12'd3001 : tab2 = 23'b10011000000110110000001;
12'd3002 : tab2 = 23'b10010111111001101101001;
12'd3003 : tab2 = 23'b10010111101100101010011;
12'd3004 : tab2 = 23'b10010111011111101000111;
12'd3005 : tab2 = 23'b10010111010010100111101;
12'd3006 : tab2 = 23'b10010111000101100111111;
12'd3007 : tab2 = 23'b10010110111000101000001;
12'd3008 : tab2 = 23'b10010110101011101000111;
12'd3009 : tab2 = 23'b10010110011110101010111;
12'd3010 : tab2 = 23'b10010110010001101101001;
12'd3011 : tab2 = 23'b10010110000100110000110;
12'd3012 : tab2 = 23'b10010101110111110100100;
12'd3013 : tab2 = 23'b10010101101010111001010;
12'd3014 : tab2 = 23'b10010101011101111110001;
12'd3015 : tab2 = 23'b10010101010001000100110;
12'd3016 : tab2 = 23'b10010101000100001011001;
12'd3017 : tab2 = 23'b10010100110111010010011;
12'd3018 : tab2 = 23'b10010100101010011010100;
12'd3019 : tab2 = 23'b10010100011101100011001;
12'd3020 : tab2 = 23'b10010100010000101100011;
12'd3021 : tab2 = 23'b10010100000011110110101;
12'd3022 : tab2 = 23'b10010011110111000001011;
12'd3023 : tab2 = 23'b10010011101010001100110;
12'd3024 : tab2 = 23'b10010011011101011000011;
12'd3025 : tab2 = 23'b10010011010000100101011;
12'd3026 : tab2 = 23'b10010011000011110010101;
12'd3027 : tab2 = 23'b10010010110111000000101;
12'd3028 : tab2 = 23'b10010010101010001111011;
12'd3029 : tab2 = 23'b10010010011101011111100;
12'd3030 : tab2 = 23'b10010010010000101111011;
12'd3031 : tab2 = 23'b10010010000011111111111;
12'd3032 : tab2 = 23'b10010001110111010001110;
12'd3033 : tab2 = 23'b10010001101010100011100;
12'd3034 : tab2 = 23'b10010001011101110110011;
12'd3035 : tab2 = 23'b10010001010001001001110;
12'd3036 : tab2 = 23'b10010001000100011110001;
12'd3037 : tab2 = 23'b10010000110111110010111;
12'd3038 : tab2 = 23'b10010000101011000111111;
12'd3039 : tab2 = 23'b10010000011110011110001;
12'd3040 : tab2 = 23'b10010000010001110101010;
12'd3041 : tab2 = 23'b10010000000101001100101;
12'd3042 : tab2 = 23'b10001111111000100100110;
12'd3043 : tab2 = 23'b10001111101011111101101;
12'd3044 : tab2 = 23'b10001111011111010110110;
12'd3045 : tab2 = 23'b10001111010010110001110;
12'd3046 : tab2 = 23'b10001111000110001100011;
12'd3047 : tab2 = 23'b10001110111001100111011;
12'd3048 : tab2 = 23'b10001110101101000100000;
12'd3049 : tab2 = 23'b10001110100000100000100;
12'd3050 : tab2 = 23'b10001110010011111101111;
12'd3051 : tab2 = 23'b10001110000111011011110;
12'd3052 : tab2 = 23'b10001101111010111010100;
12'd3053 : tab2 = 23'b10001101101110011010001;
12'd3054 : tab2 = 23'b10001101100001111010000;
12'd3055 : tab2 = 23'b10001101010101011011000;
12'd3056 : tab2 = 23'b10001101001000111100011;
12'd3057 : tab2 = 23'b10001100111100011110011;
12'd3058 : tab2 = 23'b10001100110000000000111;
12'd3059 : tab2 = 23'b10001100100011100100100;
12'd3060 : tab2 = 23'b10001100010111001000011;
12'd3061 : tab2 = 23'b10001100001010101101000;
12'd3062 : tab2 = 23'b10001011111110010001111;
12'd3063 : tab2 = 23'b10001011110001111000001;
12'd3064 : tab2 = 23'b10001011100101011110100;
12'd3065 : tab2 = 23'b10001011011001000101110;
12'd3066 : tab2 = 23'b10001011001100101110001;
12'd3067 : tab2 = 23'b10001011000000010110011;
12'd3068 : tab2 = 23'b10001010110011111111011;
12'd3069 : tab2 = 23'b10001010100111101001000;
12'd3070 : tab2 = 23'b10001010011011010011101;
12'd3071 : tab2 = 23'b10001010001110111110010;
12'd3072 : tab2 = 23'b10001010000010101010011;
12'd3073 : tab2 = 23'b10001001110110010110101;
12'd3074 : tab2 = 23'b10001001101010000100001;
12'd3075 : tab2 = 23'b10001001011101110001011;
12'd3076 : tab2 = 23'b10001001010001011111111;
12'd3077 : tab2 = 23'b10001001000101001110101;
12'd3078 : tab2 = 23'b10001000111000111110110;
12'd3079 : tab2 = 23'b10001000101100101110011;
12'd3080 : tab2 = 23'b10001000100000011111000;
12'd3081 : tab2 = 23'b10001000010100010000111;
12'd3082 : tab2 = 23'b10001000001000000010110;
12'd3083 : tab2 = 23'b10000111111011110101110;
12'd3084 : tab2 = 23'b10000111101111101000101;
12'd3085 : tab2 = 23'b10000111100011011101000;
12'd3086 : tab2 = 23'b10000111010111010001100;
12'd3087 : tab2 = 23'b10000111001011000110111;
12'd3088 : tab2 = 23'b10000110111110111100111;
12'd3089 : tab2 = 23'b10000110110010110011001;
12'd3090 : tab2 = 23'b10000110100110101010010;
12'd3091 : tab2 = 23'b10000110011010100010100;
12'd3092 : tab2 = 23'b10000110001110011010101;
12'd3093 : tab2 = 23'b10000110000010010011111;
12'd3094 : tab2 = 23'b10000101110110001101100;
12'd3095 : tab2 = 23'b10000101101010000111110;
12'd3096 : tab2 = 23'b10000101011110000010010;
12'd3097 : tab2 = 23'b10000101010001111101101;
12'd3098 : tab2 = 23'b10000101000101111010000;
12'd3099 : tab2 = 23'b10000100111001110110111;
12'd3100 : tab2 = 23'b10000100101101110100000;
12'd3101 : tab2 = 23'b10000100100001110010010;
12'd3102 : tab2 = 23'b10000100010101110000101;
12'd3103 : tab2 = 23'b10000100001001110000100;
12'd3104 : tab2 = 23'b10000011111101110000000;
12'd3105 : tab2 = 23'b10000011110001110000101;
12'd3106 : tab2 = 23'b10000011100101110001101;
12'd3107 : tab2 = 23'b10000011011001110011111;
12'd3108 : tab2 = 23'b10000011001101110101111;
12'd3109 : tab2 = 23'b10000011000001111001000;
12'd3110 : tab2 = 23'b10000010110101111100100;
12'd3111 : tab2 = 23'b10000010101010000000110;
12'd3112 : tab2 = 23'b10000010011110000101101;
12'd3113 : tab2 = 23'b10000010010010001010111;
12'd3114 : tab2 = 23'b10000010000110010000110;
12'd3115 : tab2 = 23'b10000001111010010111011;
12'd3116 : tab2 = 23'b10000001101110011110110;
12'd3117 : tab2 = 23'b10000001100010100110100;
12'd3118 : tab2 = 23'b10000001010110101110111;
12'd3119 : tab2 = 23'b10000001001010111000011;
12'd3120 : tab2 = 23'b10000000111111000001110;
12'd3121 : tab2 = 23'b10000000110011001100011;
12'd3122 : tab2 = 23'b10000000100111010111001;
12'd3123 : tab2 = 23'b10000000011011100010110;
12'd3124 : tab2 = 23'b10000000001111101111001;
12'd3125 : tab2 = 23'b10000000000011111011100;
12'd3126 : tab2 = 23'b01111111111000001000111;
12'd3127 : tab2 = 23'b01111111101100010110111;
12'd3128 : tab2 = 23'b01111111100000100101100;
12'd3129 : tab2 = 23'b01111111010100110100100;
12'd3130 : tab2 = 23'b01111111001001000100010;
12'd3131 : tab2 = 23'b01111110111101010100101;
12'd3132 : tab2 = 23'b01111110110001100101010;
12'd3133 : tab2 = 23'b01111110100101110110110;
12'd3134 : tab2 = 23'b01111110011010001000111;
12'd3135 : tab2 = 23'b01111110001110011100010;
12'd3136 : tab2 = 23'b01111110000010101111011;
12'd3137 : tab2 = 23'b01111101110111000011010;
12'd3138 : tab2 = 23'b01111101101011010111110;
12'd3139 : tab2 = 23'b01111101011111101100100;
12'd3140 : tab2 = 23'b01111101010100000010101;
12'd3141 : tab2 = 23'b01111101001000011000111;
12'd3142 : tab2 = 23'b01111100111100101111010;
12'd3143 : tab2 = 23'b01111100110001000111011;
12'd3144 : tab2 = 23'b01111100100101011110111;
12'd3145 : tab2 = 23'b01111100011001110111101;
12'd3146 : tab2 = 23'b01111100001110010001100;
12'd3147 : tab2 = 23'b01111100000010101011000;
12'd3148 : tab2 = 23'b01111011110111000110000;
12'd3149 : tab2 = 23'b01111011101011100000100;
12'd3150 : tab2 = 23'b01111011011111111100011;
12'd3151 : tab2 = 23'b01111011010100011000010;
12'd3152 : tab2 = 23'b01111011001000110101001;
12'd3153 : tab2 = 23'b01111010111101010010101;
12'd3154 : tab2 = 23'b01111010110001110000110;
12'd3155 : tab2 = 23'b01111010100110001110101;
12'd3156 : tab2 = 23'b01111010011010101101111;
12'd3157 : tab2 = 23'b01111010001111001110001;
12'd3158 : tab2 = 23'b01111010000011101101111;
12'd3159 : tab2 = 23'b01111001111000001110101;
12'd3160 : tab2 = 23'b01111001101100110000101;
12'd3161 : tab2 = 23'b01111001100001010010011;
12'd3162 : tab2 = 23'b01111001010101110101011;
12'd3163 : tab2 = 23'b01111001001010011000001;
12'd3164 : tab2 = 23'b01111000111110111100001;
12'd3165 : tab2 = 23'b01111000110011100000101;
12'd3166 : tab2 = 23'b01111000101000000101101;
12'd3167 : tab2 = 23'b01111000011100101011001;
12'd3168 : tab2 = 23'b01111000010001010001000;
12'd3169 : tab2 = 23'b01111000000101111000000;
12'd3170 : tab2 = 23'b01110111111010011111010;
12'd3171 : tab2 = 23'b01110111101111000110110;
12'd3172 : tab2 = 23'b01110111100011101111011;
12'd3173 : tab2 = 23'b01110111011000011000010;
12'd3174 : tab2 = 23'b01110111001101000001100;
12'd3175 : tab2 = 23'b01110111000001101011110;
12'd3176 : tab2 = 23'b01110110110110010110010;
12'd3177 : tab2 = 23'b01110110101011000001100;
12'd3178 : tab2 = 23'b01110110011111101101101;
12'd3179 : tab2 = 23'b01110110010100011010010;
12'd3180 : tab2 = 23'b01110110001001000110101;
12'd3181 : tab2 = 23'b01110101111101110100011;
12'd3182 : tab2 = 23'b01110101110010100010001;
12'd3183 : tab2 = 23'b01110101100111010001010;
12'd3184 : tab2 = 23'b01110101011100000000100;
12'd3185 : tab2 = 23'b01110101010000110000000;
12'd3186 : tab2 = 23'b01110101000101100000110;
12'd3187 : tab2 = 23'b01110100111010010001101;
12'd3188 : tab2 = 23'b01110100101111000010111;
12'd3189 : tab2 = 23'b01110100100011110101000;
12'd3190 : tab2 = 23'b01110100011000100111110;
12'd3191 : tab2 = 23'b01110100001101011011000;
12'd3192 : tab2 = 23'b01110100000010001110011;
12'd3193 : tab2 = 23'b01110011110111000010101;
12'd3194 : tab2 = 23'b01110011101011111000000;
12'd3195 : tab2 = 23'b01110011100000101101001;
12'd3196 : tab2 = 23'b01110011010101100011011;
12'd3197 : tab2 = 23'b01110011001010011001011;
12'd3198 : tab2 = 23'b01110010111111010000101;
12'd3199 : tab2 = 23'b01110010110100001000001;
12'd3200 : tab2 = 23'b01110010101001000000111;
12'd3201 : tab2 = 23'b01110010011101111001001;
12'd3202 : tab2 = 23'b01110010010010110010110;
12'd3203 : tab2 = 23'b01110010000111101100100;
12'd3204 : tab2 = 23'b01110001111100100111000;
12'd3205 : tab2 = 23'b01110001110001100010010;
12'd3206 : tab2 = 23'b01110001100110011101001;
12'd3207 : tab2 = 23'b01110001011011011001010;
12'd3208 : tab2 = 23'b01110001010000010110001;
12'd3209 : tab2 = 23'b01110001000101010011000;
12'd3210 : tab2 = 23'b01110000111010010000111;
12'd3211 : tab2 = 23'b01110000101111001111010;
12'd3212 : tab2 = 23'b01110000100100001101111;
12'd3213 : tab2 = 23'b01110000011001001101010;
12'd3214 : tab2 = 23'b01110000001110001101110;
12'd3215 : tab2 = 23'b01110000000011001110000;
12'd3216 : tab2 = 23'b01101111111000001110100;
12'd3217 : tab2 = 23'b01101111101101010000101;
12'd3218 : tab2 = 23'b01101111100010010010111;
12'd3219 : tab2 = 23'b01101111010111010101100;
12'd3220 : tab2 = 23'b01101111001100011000010;
12'd3221 : tab2 = 23'b01101111000001011100010;
12'd3222 : tab2 = 23'b01101110110110100000100;
12'd3223 : tab2 = 23'b01101110101011100101010;
12'd3224 : tab2 = 23'b01101110100000101010111;
12'd3225 : tab2 = 23'b01101110010101110000101;
12'd3226 : tab2 = 23'b01101110001010110111001;
12'd3227 : tab2 = 23'b01101101111111111110010;
12'd3228 : tab2 = 23'b01101101110101000101101;
12'd3229 : tab2 = 23'b01101101101010001101101;
12'd3230 : tab2 = 23'b01101101011111010110011;
12'd3231 : tab2 = 23'b01101101010100011111011;
12'd3232 : tab2 = 23'b01101101001001101001001;
12'd3233 : tab2 = 23'b01101100111110110011011;
12'd3234 : tab2 = 23'b01101100110011111110000;
12'd3235 : tab2 = 23'b01101100101001001001110;
12'd3236 : tab2 = 23'b01101100011110010101010;
12'd3237 : tab2 = 23'b01101100010011100001111;
12'd3238 : tab2 = 23'b01101100001000101110010;
12'd3239 : tab2 = 23'b01101011111101111011111;
12'd3240 : tab2 = 23'b01101011110011001010100;
12'd3241 : tab2 = 23'b01101011101000011000011;
12'd3242 : tab2 = 23'b01101011011101100111101;
12'd3243 : tab2 = 23'b01101011010010110110110;
12'd3244 : tab2 = 23'b01101011001000000111011;
12'd3245 : tab2 = 23'b01101010111101011000001;
12'd3246 : tab2 = 23'b01101010110010101001000;
12'd3247 : tab2 = 23'b01101010100111111010101;
12'd3248 : tab2 = 23'b01101010011101001101011;
12'd3249 : tab2 = 23'b01101010010010011111111;
12'd3250 : tab2 = 23'b01101010000111110010100;
12'd3251 : tab2 = 23'b01101001111101000110011;
12'd3252 : tab2 = 23'b01101001110010011010100;
12'd3253 : tab2 = 23'b01101001100111101111110;
12'd3254 : tab2 = 23'b01101001011101000101001;
12'd3255 : tab2 = 23'b01101001010010011010110;
12'd3256 : tab2 = 23'b01101001000111110001101;
12'd3257 : tab2 = 23'b01101000111101001000101;
12'd3258 : tab2 = 23'b01101000110010011111111;
12'd3259 : tab2 = 23'b01101000100111111000010;
12'd3260 : tab2 = 23'b01101000011101010000110;
12'd3261 : tab2 = 23'b01101000010010101001101;
12'd3262 : tab2 = 23'b01101000001000000011001;
12'd3263 : tab2 = 23'b01100111111101011100110;
12'd3264 : tab2 = 23'b01100111110010111000000;
12'd3265 : tab2 = 23'b01100111101000010010100;
12'd3266 : tab2 = 23'b01100111011101101110010;
12'd3267 : tab2 = 23'b01100111010011001010010;
12'd3268 : tab2 = 23'b01100111001000100111010;
12'd3269 : tab2 = 23'b01100110111110000100100;
12'd3270 : tab2 = 23'b01100110110011100001111;
12'd3271 : tab2 = 23'b01100110101001000000001;
12'd3272 : tab2 = 23'b01100110011110011111000;
12'd3273 : tab2 = 23'b01100110010011111110100;
12'd3274 : tab2 = 23'b01100110001001011101110;
12'd3275 : tab2 = 23'b01100101111110111110001;
12'd3276 : tab2 = 23'b01100101110100011110110;
12'd3277 : tab2 = 23'b01100101101010000000011;
12'd3278 : tab2 = 23'b01100101011111100010011;
12'd3279 : tab2 = 23'b01100101010101000100100;
12'd3280 : tab2 = 23'b01100101001010100110111;
12'd3281 : tab2 = 23'b01100101000000001010011;
12'd3282 : tab2 = 23'b01100100110101101110000;
12'd3283 : tab2 = 23'b01100100101011010010110;
12'd3284 : tab2 = 23'b01100100100000110111011;
12'd3285 : tab2 = 23'b01100100010110011101001;
12'd3286 : tab2 = 23'b01100100001100000010100;
12'd3287 : tab2 = 23'b01100100000001101001000;
12'd3288 : tab2 = 23'b01100011110111001111110;
12'd3289 : tab2 = 23'b01100011101100110111010;
12'd3290 : tab2 = 23'b01100011100010011111000;
12'd3291 : tab2 = 23'b01100011011000000111010;
12'd3292 : tab2 = 23'b01100011001101110000101;
12'd3293 : tab2 = 23'b01100011000011011010000;
12'd3294 : tab2 = 23'b01100010111001000100010;
12'd3295 : tab2 = 23'b01100010101110101110001;
12'd3296 : tab2 = 23'b01100010100100011001000;
12'd3297 : tab2 = 23'b01100010011010000100011;
12'd3298 : tab2 = 23'b01100010001111110000011;
12'd3299 : tab2 = 23'b01100010000101011101001;
12'd3300 : tab2 = 23'b01100001111011001010001;
12'd3301 : tab2 = 23'b01100001110000110111001;
12'd3302 : tab2 = 23'b01100001100110100100111;
12'd3303 : tab2 = 23'b01100001011100010011011;
12'd3304 : tab2 = 23'b01100001010010000010100;
12'd3305 : tab2 = 23'b01100001000111110001110;
12'd3306 : tab2 = 23'b01100000111101100001110;
12'd3307 : tab2 = 23'b01100000110011010001111;
12'd3308 : tab2 = 23'b01100000101001000010110;
12'd3309 : tab2 = 23'b01100000011110110100010;
12'd3310 : tab2 = 23'b01100000010100100101111;
12'd3311 : tab2 = 23'b01100000001010011000010;
12'd3312 : tab2 = 23'b01100000000000001011010;
12'd3313 : tab2 = 23'b01011111110101111111000;
12'd3314 : tab2 = 23'b01011111101011110010011;
12'd3315 : tab2 = 23'b01011111100001100110111;
12'd3316 : tab2 = 23'b01011111010111011011101;
12'd3317 : tab2 = 23'b01011111001101010001000;
12'd3318 : tab2 = 23'b01011111000011000110101;
12'd3319 : tab2 = 23'b01011110111000111100111;
12'd3320 : tab2 = 23'b01011110101110110100010;
12'd3321 : tab2 = 23'b01011110100100101011011;
12'd3322 : tab2 = 23'b01011110011010100010101;
12'd3323 : tab2 = 23'b01011110010000011011101;
12'd3324 : tab2 = 23'b01011110000110010100001;
12'd3325 : tab2 = 23'b01011101111100001101011;
12'd3326 : tab2 = 23'b01011101110010000111010;
12'd3327 : tab2 = 23'b01011101101000000001000;
12'd3328 : tab2 = 23'b01011101011101111011110;
12'd3329 : tab2 = 23'b01011101010011110110101;
12'd3330 : tab2 = 23'b01011101001001110010110;
12'd3331 : tab2 = 23'b01011100111111101111001;
12'd3332 : tab2 = 23'b01011100110101101011100;
12'd3333 : tab2 = 23'b01011100101011101000001;
12'd3334 : tab2 = 23'b01011100100001100110000;
12'd3335 : tab2 = 23'b01011100010111100011111;
12'd3336 : tab2 = 23'b01011100001101100010100;
12'd3337 : tab2 = 23'b01011100000011100001111;
12'd3338 : tab2 = 23'b01011011111001100000110;
12'd3339 : tab2 = 23'b01011011101111100001010;
12'd3340 : tab2 = 23'b01011011100101100001110;
12'd3341 : tab2 = 23'b01011011011011100010101;
12'd3342 : tab2 = 23'b01011011010001100100010;
12'd3343 : tab2 = 23'b01011011000111100110000;
12'd3344 : tab2 = 23'b01011010111101101000100;
12'd3345 : tab2 = 23'b01011010110011101011001;
12'd3346 : tab2 = 23'b01011010101001101110100;
12'd3347 : tab2 = 23'b01011010011111110010011;
12'd3348 : tab2 = 23'b01011010010101110110100;
12'd3349 : tab2 = 23'b01011010001011111011010;
12'd3350 : tab2 = 23'b01011010000010000000110;
12'd3351 : tab2 = 23'b01011001111000000110011;
12'd3352 : tab2 = 23'b01011001101110001100100;
12'd3353 : tab2 = 23'b01011001100100010011000;
12'd3354 : tab2 = 23'b01011001011010011010101;
12'd3355 : tab2 = 23'b01011001010000100001111;
12'd3356 : tab2 = 23'b01011001000110101001110;
12'd3357 : tab2 = 23'b01011000111100110010011;
12'd3358 : tab2 = 23'b01011000110010111011101;
12'd3359 : tab2 = 23'b01011000101001000101000;
12'd3360 : tab2 = 23'b01011000011111001110101;
12'd3361 : tab2 = 23'b01011000010101011000110;
12'd3362 : tab2 = 23'b01011000001011100100010;
12'd3363 : tab2 = 23'b01011000000001101111110;
12'd3364 : tab2 = 23'b01010111110111111011100;
12'd3365 : tab2 = 23'b01010111101110000111011;
12'd3366 : tab2 = 23'b01010111100100010100010;
12'd3367 : tab2 = 23'b01010111011010100001100;
12'd3368 : tab2 = 23'b01010111010000101110111;
12'd3369 : tab2 = 23'b01010111000110111101011;
12'd3370 : tab2 = 23'b01010110111101001100000;
12'd3371 : tab2 = 23'b01010110110011011010111;
12'd3372 : tab2 = 23'b01010110101001101010011;
12'd3373 : tab2 = 23'b01010110011111111010100;
12'd3374 : tab2 = 23'b01010110010110001010111;
12'd3375 : tab2 = 23'b01010110001100011011111;
12'd3376 : tab2 = 23'b01010110000010101101011;
12'd3377 : tab2 = 23'b01010101111000111111001;
12'd3378 : tab2 = 23'b01010101101111010001001;
12'd3379 : tab2 = 23'b01010101100101100100001;
12'd3380 : tab2 = 23'b01010101011011110111100;
12'd3381 : tab2 = 23'b01010101010010001010111;
12'd3382 : tab2 = 23'b01010101001000011111010;
12'd3383 : tab2 = 23'b01010100111110110011101;
12'd3384 : tab2 = 23'b01010100110101001000111;
12'd3385 : tab2 = 23'b01010100101011011110100;
12'd3386 : tab2 = 23'b01010100100001110100010;
12'd3387 : tab2 = 23'b01010100011000001010100;
12'd3388 : tab2 = 23'b01010100001110100001111;
12'd3389 : tab2 = 23'b01010100000100111000101;
12'd3390 : tab2 = 23'b01010011111011010000011;
12'd3391 : tab2 = 23'b01010011110001101001010;
12'd3392 : tab2 = 23'b01010011101000000001100;
12'd3393 : tab2 = 23'b01010011011110011010110;
12'd3394 : tab2 = 23'b01010011010100110100001;
12'd3395 : tab2 = 23'b01010011001011001110101;
12'd3396 : tab2 = 23'b01010011000001101000110;
12'd3397 : tab2 = 23'b01010010111000000011101;
12'd3398 : tab2 = 23'b01010010101110011111001;
12'd3399 : tab2 = 23'b01010010100100111011010;
12'd3400 : tab2 = 23'b01010010011011010111101;
12'd3401 : tab2 = 23'b01010010010001110100001;
12'd3402 : tab2 = 23'b01010010001000010001010;
12'd3403 : tab2 = 23'b01010001111110101110111;
12'd3404 : tab2 = 23'b01010001110101001101011;
12'd3405 : tab2 = 23'b01010001101011101011100;
12'd3406 : tab2 = 23'b01010001100010001010101;
12'd3407 : tab2 = 23'b01010001011000101010001;
12'd3408 : tab2 = 23'b01010001001111001010001;
12'd3409 : tab2 = 23'b01010001000101101010001;
12'd3410 : tab2 = 23'b01010000111100001011001;
12'd3411 : tab2 = 23'b01010000110010101100000;
12'd3412 : tab2 = 23'b01010000101001001110001;
12'd3413 : tab2 = 23'b01010000011111110000011;
12'd3414 : tab2 = 23'b01010000010110010010110;
12'd3415 : tab2 = 23'b01010000001100110101011;
12'd3416 : tab2 = 23'b01010000000011011001000;
12'd3417 : tab2 = 23'b01001111111001111100110;
12'd3418 : tab2 = 23'b01001111110000100001011;
12'd3419 : tab2 = 23'b01001111100111000110000;
12'd3420 : tab2 = 23'b01001111011101101011010;
12'd3421 : tab2 = 23'b01001111010100010000110;
12'd3422 : tab2 = 23'b01001111001010110111010;
12'd3423 : tab2 = 23'b01001111000001011101100;
12'd3424 : tab2 = 23'b01001110111000000100111;
12'd3425 : tab2 = 23'b01001110101110101011111;
12'd3426 : tab2 = 23'b01001110100101010100000;
12'd3427 : tab2 = 23'b01001110011011111100011;
12'd3428 : tab2 = 23'b01001110010010100100110;
12'd3429 : tab2 = 23'b01001110001001001101111;
12'd3430 : tab2 = 23'b01001101111111110111101;
12'd3431 : tab2 = 23'b01001101110110100010000;
12'd3432 : tab2 = 23'b01001101101101001100000;
12'd3433 : tab2 = 23'b01001101100011110111001;
12'd3434 : tab2 = 23'b01001101011010100010100;
12'd3435 : tab2 = 23'b01001101010001001101111;
12'd3436 : tab2 = 23'b01001101000111111010000;
12'd3437 : tab2 = 23'b01001100111110100110110;
12'd3438 : tab2 = 23'b01001100110101010100001;
12'd3439 : tab2 = 23'b01001100101100000001001;
12'd3440 : tab2 = 23'b01001100100010101111011;
12'd3441 : tab2 = 23'b01001100011001011101101;
12'd3442 : tab2 = 23'b01001100010000001100001;
12'd3443 : tab2 = 23'b01001100000110111011110;
12'd3444 : tab2 = 23'b01001011111101101011011;
12'd3445 : tab2 = 23'b01001011110100011011010;
12'd3446 : tab2 = 23'b01001011101011001100010;
12'd3447 : tab2 = 23'b01001011100001111101000;
12'd3448 : tab2 = 23'b01001011011000101110110;
12'd3449 : tab2 = 23'b01001011001111100000001;
12'd3450 : tab2 = 23'b01001011000110010010101;
12'd3451 : tab2 = 23'b01001010111101000101011;
12'd3452 : tab2 = 23'b01001010110011111000010;
12'd3453 : tab2 = 23'b01001010101010101011011;
12'd3454 : tab2 = 23'b01001010100001011111100;
12'd3455 : tab2 = 23'b01001010011000010011110;
12'd3456 : tab2 = 23'b01001010001111001001000;
12'd3457 : tab2 = 23'b01001010000101111110001;
12'd3458 : tab2 = 23'b01001001111100110011110;
12'd3459 : tab2 = 23'b01001001110011101010000;
12'd3460 : tab2 = 23'b01001001101010100000001;
12'd3461 : tab2 = 23'b01001001100001010111001;
12'd3462 : tab2 = 23'b01001001011000001110011;
12'd3463 : tab2 = 23'b01001001001111000101110;
12'd3464 : tab2 = 23'b01001001000101111110010;
12'd3465 : tab2 = 23'b01001000111100110110111;
12'd3466 : tab2 = 23'b01001000110011101111101;
12'd3467 : tab2 = 23'b01001000101010101001100;
12'd3468 : tab2 = 23'b01001000100001100011000;
12'd3469 : tab2 = 23'b01001000011000011101110;
12'd3470 : tab2 = 23'b01001000001111011000001;
12'd3471 : tab2 = 23'b01001000000110010011100;
12'd3472 : tab2 = 23'b01000111111101001110101;
12'd3473 : tab2 = 23'b01000111110100001010110;
12'd3474 : tab2 = 23'b01000111101011000111001;
12'd3475 : tab2 = 23'b01000111100010000011110;
12'd3476 : tab2 = 23'b01000111011001000000111;
12'd3477 : tab2 = 23'b01000111001111111110111;
12'd3478 : tab2 = 23'b01000111000110111100011;
12'd3479 : tab2 = 23'b01000110111101111011000;
12'd3480 : tab2 = 23'b01000110110100111010001;
12'd3481 : tab2 = 23'b01000110101011111001011;
12'd3482 : tab2 = 23'b01000110100010111000110;
12'd3483 : tab2 = 23'b01000110011001111001011;
12'd3484 : tab2 = 23'b01000110010000111001100;
12'd3485 : tab2 = 23'b01000110000111111010011;
12'd3486 : tab2 = 23'b01000101111110111011110;
12'd3487 : tab2 = 23'b01000101110101111101110;
12'd3488 : tab2 = 23'b01000101101100111111100;
12'd3489 : tab2 = 23'b01000101100100000010011;
12'd3490 : tab2 = 23'b01000101011011000101011;
12'd3491 : tab2 = 23'b01000101010010001000100;
12'd3492 : tab2 = 23'b01000101001001001100101;
12'd3493 : tab2 = 23'b01000101000000010000101;
12'd3494 : tab2 = 23'b01000100110111010101100;
12'd3495 : tab2 = 23'b01000100101110011010001;
12'd3496 : tab2 = 23'b01000100100101011111111;
12'd3497 : tab2 = 23'b01000100011100100101111;
12'd3498 : tab2 = 23'b01000100010011101011110;
12'd3499 : tab2 = 23'b01000100001010110010100;
12'd3500 : tab2 = 23'b01000100000001111001110;
12'd3501 : tab2 = 23'b01000011111001000000101;
12'd3502 : tab2 = 23'b01000011110000001001001;
12'd3503 : tab2 = 23'b01000011100111010001001;
12'd3504 : tab2 = 23'b01000011011110011001100;
12'd3505 : tab2 = 23'b01000011010101100011011;
12'd3506 : tab2 = 23'b01000011001100101100100;
12'd3507 : tab2 = 23'b01000011000011110110101;
12'd3508 : tab2 = 23'b01000010111011000000111;
12'd3509 : tab2 = 23'b01000010110010001011011;
12'd3510 : tab2 = 23'b01000010101001010110011;
12'd3511 : tab2 = 23'b01000010100000100010000;
12'd3512 : tab2 = 23'b01000010010111101110010;
12'd3513 : tab2 = 23'b01000010001110111010010;
12'd3514 : tab2 = 23'b01000010000110000110111;
12'd3515 : tab2 = 23'b01000001111101010100000;
12'd3516 : tab2 = 23'b01000001110100100001110;
12'd3517 : tab2 = 23'b01000001101011101111010;
12'd3518 : tab2 = 23'b01000001100010111101110;
12'd3519 : tab2 = 23'b01000001011010001100100;
12'd3520 : tab2 = 23'b01000001010001011100001;
12'd3521 : tab2 = 23'b01000001001000101011001;
12'd3522 : tab2 = 23'b01000000111111111011001;
12'd3523 : tab2 = 23'b01000000110111001011010;
12'd3524 : tab2 = 23'b01000000101110011100001;
12'd3525 : tab2 = 23'b01000000100101101101001;
12'd3526 : tab2 = 23'b01000000011100111110100;
12'd3527 : tab2 = 23'b01000000010100010000010;
12'd3528 : tab2 = 23'b01000000001011100011000;
12'd3529 : tab2 = 23'b01000000000010110101111;
12'd3530 : tab2 = 23'b00111111111010001000111;
12'd3531 : tab2 = 23'b00111111110001011100001;
12'd3532 : tab2 = 23'b00111111101000101111111;
12'd3533 : tab2 = 23'b00111111100000000100010;
12'd3534 : tab2 = 23'b00111111010111011001010;
12'd3535 : tab2 = 23'b00111111001110101101111;
12'd3536 : tab2 = 23'b00111111000110000011110;
12'd3537 : tab2 = 23'b00111110111101011001100;
12'd3538 : tab2 = 23'b00111110110100101111100;
12'd3539 : tab2 = 23'b00111110101100000101110;
12'd3540 : tab2 = 23'b00111110100011011101000;
12'd3541 : tab2 = 23'b00111110011010110100011;
12'd3542 : tab2 = 23'b00111110010010001100011;
12'd3543 : tab2 = 23'b00111110001001100100011;
12'd3544 : tab2 = 23'b00111110000000111101001;
12'd3545 : tab2 = 23'b00111101111000010110000;
12'd3546 : tab2 = 23'b00111101101111101111000;
12'd3547 : tab2 = 23'b00111101100111001001000;
12'd3548 : tab2 = 23'b00111101011110100011010;
12'd3549 : tab2 = 23'b00111101010101111101100;
12'd3550 : tab2 = 23'b00111101001101011000001;
12'd3551 : tab2 = 23'b00111101000100110011100;
12'd3552 : tab2 = 23'b00111100111100001111010;
12'd3553 : tab2 = 23'b00111100110011101011001;
12'd3554 : tab2 = 23'b00111100101011001000000;
12'd3555 : tab2 = 23'b00111100100010100101000;
12'd3556 : tab2 = 23'b00111100011010000010001;
12'd3557 : tab2 = 23'b00111100010001011111011;
12'd3558 : tab2 = 23'b00111100001000111101110;
12'd3559 : tab2 = 23'b00111100000000011011110;
12'd3560 : tab2 = 23'b00111011110111111010110;
12'd3561 : tab2 = 23'b00111011101111011001101;
12'd3562 : tab2 = 23'b00111011100110111001000;
12'd3563 : tab2 = 23'b00111011011110011001000;
12'd3564 : tab2 = 23'b00111011010101111001101;
12'd3565 : tab2 = 23'b00111011001101011001110;
12'd3566 : tab2 = 23'b00111011000100111011000;
12'd3567 : tab2 = 23'b00111010111100011100100;
12'd3568 : tab2 = 23'b00111010110011111110001;
12'd3569 : tab2 = 23'b00111010101011100000110;
12'd3570 : tab2 = 23'b00111010100011000010111;
12'd3571 : tab2 = 23'b00111010011010100101111;
12'd3572 : tab2 = 23'b00111010010010001001011;
12'd3573 : tab2 = 23'b00111010001001101100100;
12'd3574 : tab2 = 23'b00111010000001010000110;
12'd3575 : tab2 = 23'b00111001111000110101001;
12'd3576 : tab2 = 23'b00111001110000011010001;
12'd3577 : tab2 = 23'b00111001100111111111001;
12'd3578 : tab2 = 23'b00111001011111100100110;
12'd3579 : tab2 = 23'b00111001010111001010101;
12'd3580 : tab2 = 23'b00111001001110110001100;
12'd3581 : tab2 = 23'b00111001000110010111100;
12'd3582 : tab2 = 23'b00111000111101111110110;
12'd3583 : tab2 = 23'b00111000110101100110100;
12'd3584 : tab2 = 23'b00111000101101001110010;
12'd3585 : tab2 = 23'b00111000100100110110011;
12'd3586 : tab2 = 23'b00111000011100011110111;
12'd3587 : tab2 = 23'b00111000010100001000000;
12'd3588 : tab2 = 23'b00111000001011110001010;
12'd3589 : tab2 = 23'b00111000000011011010111;
12'd3590 : tab2 = 23'b00110111111011000100111;
12'd3591 : tab2 = 23'b00110111110010101111011;
12'd3592 : tab2 = 23'b00110111101010011010010;
12'd3593 : tab2 = 23'b00110111100010000101100;
12'd3594 : tab2 = 23'b00110111011001110001000;
12'd3595 : tab2 = 23'b00110111010001011100101;
12'd3596 : tab2 = 23'b00110111001001001001010;
12'd3597 : tab2 = 23'b00110111000000110101101;
12'd3598 : tab2 = 23'b00110110111000100011000;
12'd3599 : tab2 = 23'b00110110110000010000001;
12'd3600 : tab2 = 23'b00110110100111111110001;
12'd3601 : tab2 = 23'b00110110011111101100000;
12'd3602 : tab2 = 23'b00110110010111011010110;
12'd3603 : tab2 = 23'b00110110001111001001010;
12'd3604 : tab2 = 23'b00110110000110111000111;
12'd3605 : tab2 = 23'b00110101111110101000100;
12'd3606 : tab2 = 23'b00110101110110011000010;
12'd3607 : tab2 = 23'b00110101101110001000010;
12'd3608 : tab2 = 23'b00110101100101111001010;
12'd3609 : tab2 = 23'b00110101011101101010010;
12'd3610 : tab2 = 23'b00110101010101011011101;
12'd3611 : tab2 = 23'b00110101001101001101011;
12'd3612 : tab2 = 23'b00110101000100111111010;
12'd3613 : tab2 = 23'b00110100111100110010010;
12'd3614 : tab2 = 23'b00110100110100100101000;
12'd3615 : tab2 = 23'b00110100101100011000010;
12'd3616 : tab2 = 23'b00110100100100001011101;
12'd3617 : tab2 = 23'b00110100011100000000001;
12'd3618 : tab2 = 23'b00110100010011110100010;
12'd3619 : tab2 = 23'b00110100001011101000111;
12'd3620 : tab2 = 23'b00110100000011011110001;
12'd3621 : tab2 = 23'b00110011111011010011011;
12'd3622 : tab2 = 23'b00110011110011001001000;
12'd3623 : tab2 = 23'b00110011101010111111001;
12'd3624 : tab2 = 23'b00110011100010110101110;
12'd3625 : tab2 = 23'b00110011011010101100101;
12'd3626 : tab2 = 23'b00110011010010100011101;
12'd3627 : tab2 = 23'b00110011001010011011101;
12'd3628 : tab2 = 23'b00110011000010010011010;
12'd3629 : tab2 = 23'b00110010111010001011100;
12'd3630 : tab2 = 23'b00110010110010000100010;
12'd3631 : tab2 = 23'b00110010101001111101001;
12'd3632 : tab2 = 23'b00110010100001110110010;
12'd3633 : tab2 = 23'b00110010011001110000000;
12'd3634 : tab2 = 23'b00110010010001101010101;
12'd3635 : tab2 = 23'b00110010001001100100100;
12'd3636 : tab2 = 23'b00110010000001011111100;
12'd3637 : tab2 = 23'b00110001111001011010100;
12'd3638 : tab2 = 23'b00110001110001010110010;
12'd3639 : tab2 = 23'b00110001101001010001111;
12'd3640 : tab2 = 23'b00110001100001001110011;
12'd3641 : tab2 = 23'b00110001011001001010111;
12'd3642 : tab2 = 23'b00110001010001000111011;
12'd3643 : tab2 = 23'b00110001001001000101001;
12'd3644 : tab2 = 23'b00110001000001000010111;
12'd3645 : tab2 = 23'b00110000111001000000101;
12'd3646 : tab2 = 23'b00110000110000111110110;
12'd3647 : tab2 = 23'b00110000101000111101101;
12'd3648 : tab2 = 23'b00110000100000111100100;
12'd3649 : tab2 = 23'b00110000011000111100001;
12'd3650 : tab2 = 23'b00110000010000111011101;
12'd3651 : tab2 = 23'b00110000001000111100001;
12'd3652 : tab2 = 23'b00110000000000111100001;
12'd3653 : tab2 = 23'b00101111111000111101011;
12'd3654 : tab2 = 23'b00101111110000111110001;
12'd3655 : tab2 = 23'b00101111101000111111101;
12'd3656 : tab2 = 23'b00101111100001000001100;
12'd3657 : tab2 = 23'b00101111011001000011101;
12'd3658 : tab2 = 23'b00101111010001000110010;
12'd3659 : tab2 = 23'b00101111001001001001000;
12'd3660 : tab2 = 23'b00101111000001001100100;
12'd3661 : tab2 = 23'b00101110111001001111100;
12'd3662 : tab2 = 23'b00101110110001010011111;
12'd3663 : tab2 = 23'b00101110101001010111110;
12'd3664 : tab2 = 23'b00101110100001011100100;
12'd3665 : tab2 = 23'b00101110011001100001011;
12'd3666 : tab2 = 23'b00101110010001100111010;
12'd3667 : tab2 = 23'b00101110001001101100100;
12'd3668 : tab2 = 23'b00101110000001110010100;
12'd3669 : tab2 = 23'b00101101111001111000111;
12'd3670 : tab2 = 23'b00101101110001111111010;
12'd3671 : tab2 = 23'b00101101101010000110110;
12'd3672 : tab2 = 23'b00101101100010001101110;
12'd3673 : tab2 = 23'b00101101011010010101111;
12'd3674 : tab2 = 23'b00101101010010011101101;
12'd3675 : tab2 = 23'b00101101001010100110011;
12'd3676 : tab2 = 23'b00101101000010101110111;
12'd3677 : tab2 = 23'b00101100111010111000000;
12'd3678 : tab2 = 23'b00101100110011000001101;
12'd3679 : tab2 = 23'b00101100101011001010111;
12'd3680 : tab2 = 23'b00101100100011010101010;
12'd3681 : tab2 = 23'b00101100011011011111101;
12'd3682 : tab2 = 23'b00101100010011101010001;
12'd3683 : tab2 = 23'b00101100001011110101110;
12'd3684 : tab2 = 23'b00101100000100000001000;
12'd3685 : tab2 = 23'b00101011111100001100110;
12'd3686 : tab2 = 23'b00101011110100011001001;
12'd3687 : tab2 = 23'b00101011101100100101010;
12'd3688 : tab2 = 23'b00101011100100110010011;
12'd3689 : tab2 = 23'b00101011011100111111100;
12'd3690 : tab2 = 23'b00101011010101001100110;
12'd3691 : tab2 = 23'b00101011001101011010110;
12'd3692 : tab2 = 23'b00101011000101101000101;
12'd3693 : tab2 = 23'b00101010111101110111010;
12'd3694 : tab2 = 23'b00101010110110000101111;
12'd3695 : tab2 = 23'b00101010101110010101101;
12'd3696 : tab2 = 23'b00101010100110100101000;
12'd3697 : tab2 = 23'b00101010011110110100111;
12'd3698 : tab2 = 23'b00101010010111000101000;
12'd3699 : tab2 = 23'b00101010001111010101100;
12'd3700 : tab2 = 23'b00101010000111100110011;
12'd3701 : tab2 = 23'b00101001111111110111101;
12'd3702 : tab2 = 23'b00101001111000001001011;
12'd3703 : tab2 = 23'b00101001110000011011000;
12'd3704 : tab2 = 23'b00101001101000101101001;
12'd3705 : tab2 = 23'b00101001100000111111110;
12'd3706 : tab2 = 23'b00101001011001010011000;
12'd3707 : tab2 = 23'b00101001010001100101111;
12'd3708 : tab2 = 23'b00101001001001111001011;
12'd3709 : tab2 = 23'b00101001000010001101000;
12'd3710 : tab2 = 23'b00101000111010100001001;
12'd3711 : tab2 = 23'b00101000110010110110010;
12'd3712 : tab2 = 23'b00101000101011001010101;
12'd3713 : tab2 = 23'b00101000100011100000000;
12'd3714 : tab2 = 23'b00101000011011110101100;
12'd3715 : tab2 = 23'b00101000010100001011001;
12'd3716 : tab2 = 23'b00101000001100100001110;
12'd3717 : tab2 = 23'b00101000000100111000000;
12'd3718 : tab2 = 23'b00100111111101001110101;
12'd3719 : tab2 = 23'b00100111110101100101111;
12'd3720 : tab2 = 23'b00100111101101111101100;
12'd3721 : tab2 = 23'b00100111100110010101000;
12'd3722 : tab2 = 23'b00100111011110101101110;
12'd3723 : tab2 = 23'b00100111010111000110001;
12'd3724 : tab2 = 23'b00100111001111011110101;
12'd3725 : tab2 = 23'b00100111000111111000000;
12'd3726 : tab2 = 23'b00100111000000010001001;
12'd3727 : tab2 = 23'b00100110111000101011010;
12'd3728 : tab2 = 23'b00100110110001000101001;
12'd3729 : tab2 = 23'b00100110101001011111111;
12'd3730 : tab2 = 23'b00100110100001111010011;
12'd3731 : tab2 = 23'b00100110011010010101110;
12'd3732 : tab2 = 23'b00100110010010110000111;
12'd3733 : tab2 = 23'b00100110001011001100101;
12'd3734 : tab2 = 23'b00100110000011101000100;
12'd3735 : tab2 = 23'b00100101111100000100111;
12'd3736 : tab2 = 23'b00100101110100100010001;
12'd3737 : tab2 = 23'b00100101101100111110111;
12'd3738 : tab2 = 23'b00100101100101011100000;
12'd3739 : tab2 = 23'b00100101011101111010000;
12'd3740 : tab2 = 23'b00100101010110010111111;
12'd3741 : tab2 = 23'b00100101001110110101111;
12'd3742 : tab2 = 23'b00100101000111010100111;
12'd3743 : tab2 = 23'b00100100111111110011111;
12'd3744 : tab2 = 23'b00100100111000010011000;
12'd3745 : tab2 = 23'b00100100110000110010011;
12'd3746 : tab2 = 23'b00100100101001010010101;
12'd3747 : tab2 = 23'b00100100100001110010101;
12'd3748 : tab2 = 23'b00100100011010010011100;
12'd3749 : tab2 = 23'b00100100010010110100001;
12'd3750 : tab2 = 23'b00100100001011010101011;
12'd3751 : tab2 = 23'b00100100000011110110110;
12'd3752 : tab2 = 23'b00100011111100011000100;
12'd3753 : tab2 = 23'b00100011110100111010011;
12'd3754 : tab2 = 23'b00100011101101011101011;
12'd3755 : tab2 = 23'b00100011100110000000011;
12'd3756 : tab2 = 23'b00100011011110100011101;
12'd3757 : tab2 = 23'b00100011010111000110111;
12'd3758 : tab2 = 23'b00100011001111101010010;
12'd3759 : tab2 = 23'b00100011001000001110101;
12'd3760 : tab2 = 23'b00100011000000110010110;
12'd3761 : tab2 = 23'b00100010111001010111111;
12'd3762 : tab2 = 23'b00100010110001111100101;
12'd3763 : tab2 = 23'b00100010101010100001111;
12'd3764 : tab2 = 23'b00100010100011000111101;
12'd3765 : tab2 = 23'b00100010011011101101100;
12'd3766 : tab2 = 23'b00100010010100010100001;
12'd3767 : tab2 = 23'b00100010001100111010001;
12'd3768 : tab2 = 23'b00100010000101100001011;
12'd3769 : tab2 = 23'b00100001111110001000101;
12'd3770 : tab2 = 23'b00100001110110110000000;
12'd3771 : tab2 = 23'b00100001101111010111111;
12'd3772 : tab2 = 23'b00100001101000000000000;
12'd3773 : tab2 = 23'b00100001100000101000100;
12'd3774 : tab2 = 23'b00100001011001010001010;
12'd3775 : tab2 = 23'b00100001010001111010000;
12'd3776 : tab2 = 23'b00100001001010100011110;
12'd3777 : tab2 = 23'b00100001000011001101010;
12'd3778 : tab2 = 23'b00100000111011110111110;
12'd3779 : tab2 = 23'b00100000110100100001111;
12'd3780 : tab2 = 23'b00100000101101001100101;
12'd3781 : tab2 = 23'b00100000100101110111010;
12'd3782 : tab2 = 23'b00100000011110100010101;
12'd3783 : tab2 = 23'b00100000010111001110001;
12'd3784 : tab2 = 23'b00100000001111111010100;
12'd3785 : tab2 = 23'b00100000001000100110010;
12'd3786 : tab2 = 23'b00100000000001010010110;
12'd3787 : tab2 = 23'b00011111111001111111100;
12'd3788 : tab2 = 23'b00011111110010101100011;
12'd3789 : tab2 = 23'b00011111101011011010010;
12'd3790 : tab2 = 23'b00011111100100000111110;
12'd3791 : tab2 = 23'b00011111011100110101110;
12'd3792 : tab2 = 23'b00011111010101100100011;
12'd3793 : tab2 = 23'b00011111001110010010110;
12'd3794 : tab2 = 23'b00011111000111000001111;
12'd3795 : tab2 = 23'b00011110111111110001011;
12'd3796 : tab2 = 23'b00011110111000100000110;
12'd3797 : tab2 = 23'b00011110110001010000011;
12'd3798 : tab2 = 23'b00011110101010000000111;
12'd3799 : tab2 = 23'b00011110100010110001001;
12'd3800 : tab2 = 23'b00011110011011100010010;
12'd3801 : tab2 = 23'b00011110010100010011010;
12'd3802 : tab2 = 23'b00011110001101000100101;
12'd3803 : tab2 = 23'b00011110000101110110010;
12'd3804 : tab2 = 23'b00011101111110101000010;
12'd3805 : tab2 = 23'b00011101110111011010011;
12'd3806 : tab2 = 23'b00011101110000001101100;
12'd3807 : tab2 = 23'b00011101101001000000000;
12'd3808 : tab2 = 23'b00011101100001110011011;
12'd3809 : tab2 = 23'b00011101011010100110110;
12'd3810 : tab2 = 23'b00011101010011011010011;
12'd3811 : tab2 = 23'b00011101001100001111000;
12'd3812 : tab2 = 23'b00011101000101000011010;
12'd3813 : tab2 = 23'b00011100111101111000011;
12'd3814 : tab2 = 23'b00011100110110101101010;
12'd3815 : tab2 = 23'b00011100101111100010010;
12'd3816 : tab2 = 23'b00011100101000011000010;
12'd3817 : tab2 = 23'b00011100100001001101111;
12'd3818 : tab2 = 23'b00011100011010000100100;
12'd3819 : tab2 = 23'b00011100010010111010110;
12'd3820 : tab2 = 23'b00011100001011110001101;
12'd3821 : tab2 = 23'b00011100000100101000100;
12'd3822 : tab2 = 23'b00011011111101011111111;
12'd3823 : tab2 = 23'b00011011110110010111101;
12'd3824 : tab2 = 23'b00011011101111010000000;
12'd3825 : tab2 = 23'b00011011101000001000010;
12'd3826 : tab2 = 23'b00011011100001000001000;
12'd3827 : tab2 = 23'b00011011011001111001111;
12'd3828 : tab2 = 23'b00011011010010110011010;
12'd3829 : tab2 = 23'b00011011001011101100011;
12'd3830 : tab2 = 23'b00011011000100100110011;
12'd3831 : tab2 = 23'b00011010111101100000100;
12'd3832 : tab2 = 23'b00011010110110011010110;
12'd3833 : tab2 = 23'b00011010101111010101100;
12'd3834 : tab2 = 23'b00011010101000010000011;
12'd3835 : tab2 = 23'b00011010100001001011111;
12'd3836 : tab2 = 23'b00011010011010000111011;
12'd3837 : tab2 = 23'b00011010010011000011000;
12'd3838 : tab2 = 23'b00011010001011111111101;
12'd3839 : tab2 = 23'b00011010000100111100010;
12'd3840 : tab2 = 23'b00011001111101111001000;
12'd3841 : tab2 = 23'b00011001110110110110000;
12'd3842 : tab2 = 23'b00011001101111110011000;
12'd3843 : tab2 = 23'b00011001101000110000111;
12'd3844 : tab2 = 23'b00011001100001101111000;
12'd3845 : tab2 = 23'b00011001011010101101001;
12'd3846 : tab2 = 23'b00011001010011101011100;
12'd3847 : tab2 = 23'b00011001001100101010000;
12'd3848 : tab2 = 23'b00011001000101101001010;
12'd3849 : tab2 = 23'b00011000111110101000101;
12'd3850 : tab2 = 23'b00011000110111101000011;
12'd3851 : tab2 = 23'b00011000110000101000110;
12'd3852 : tab2 = 23'b00011000101001101000100;
12'd3853 : tab2 = 23'b00011000100010101001011;
12'd3854 : tab2 = 23'b00011000011011101010001;
12'd3855 : tab2 = 23'b00011000010100101011000;
12'd3856 : tab2 = 23'b00011000001101101100111;
12'd3857 : tab2 = 23'b00011000000110101110100;
12'd3858 : tab2 = 23'b00010111111111110000101;
12'd3859 : tab2 = 23'b00010111111000110011001;
12'd3860 : tab2 = 23'b00010111110001110101100;
12'd3861 : tab2 = 23'b00010111101010111000011;
12'd3862 : tab2 = 23'b00010111100011111011010;
12'd3863 : tab2 = 23'b00010111011100111110110;
12'd3864 : tab2 = 23'b00010111010110000010010;
12'd3865 : tab2 = 23'b00010111001111000110111;
12'd3866 : tab2 = 23'b00010111001000001011000;
12'd3867 : tab2 = 23'b00010111000001001111011;
12'd3868 : tab2 = 23'b00010110111010010100001;
12'd3869 : tab2 = 23'b00010110110011011001101;
12'd3870 : tab2 = 23'b00010110101100011110111;
12'd3871 : tab2 = 23'b00010110100101100101000;
12'd3872 : tab2 = 23'b00010110011110101011000;
12'd3873 : tab2 = 23'b00010110010111110001010;
12'd3874 : tab2 = 23'b00010110010000110111101;
12'd3875 : tab2 = 23'b00010110001001111110110;
12'd3876 : tab2 = 23'b00010110000011000101110;
12'd3877 : tab2 = 23'b00010101111100001101100;
12'd3878 : tab2 = 23'b00010101110101010101000;
12'd3879 : tab2 = 23'b00010101101110011101001;
12'd3880 : tab2 = 23'b00010101100111100101011;
12'd3881 : tab2 = 23'b00010101100000101110000;
12'd3882 : tab2 = 23'b00010101011001110110111;
12'd3883 : tab2 = 23'b00010101010010111111110;
12'd3884 : tab2 = 23'b00010101001100001001100;
12'd3885 : tab2 = 23'b00010101000101010011001;
12'd3886 : tab2 = 23'b00010100111110011101001;
12'd3887 : tab2 = 23'b00010100110111100111011;
12'd3888 : tab2 = 23'b00010100110000110010000;
12'd3889 : tab2 = 23'b00010100101001111100110;
12'd3890 : tab2 = 23'b00010100100011000111110;
12'd3891 : tab2 = 23'b00010100011100010011000;
12'd3892 : tab2 = 23'b00010100010101011111000;
12'd3893 : tab2 = 23'b00010100001110101011000;
12'd3894 : tab2 = 23'b00010100000111110111000;
12'd3895 : tab2 = 23'b00010100000001000011110;
12'd3896 : tab2 = 23'b00010011111010010000111;
12'd3897 : tab2 = 23'b00010011110011011101110;
12'd3898 : tab2 = 23'b00010011101100101010110;
12'd3899 : tab2 = 23'b00010011100101111000101;
12'd3900 : tab2 = 23'b00010011011111000110100;
12'd3901 : tab2 = 23'b00010011011000010100101;
12'd3902 : tab2 = 23'b00010011010001100011010;
12'd3903 : tab2 = 23'b00010011001010110010000;
12'd3904 : tab2 = 23'b00010011000100000000111;
12'd3905 : tab2 = 23'b00010010111101010000100;
12'd3906 : tab2 = 23'b00010010110110100000000;
12'd3907 : tab2 = 23'b00010010101111101111100;
12'd3908 : tab2 = 23'b00010010101001000000000;
12'd3909 : tab2 = 23'b00010010100010010000100;
12'd3910 : tab2 = 23'b00010010011011100001001;
12'd3911 : tab2 = 23'b00010010010100110001111;
12'd3912 : tab2 = 23'b00010010001110000011010;
12'd3913 : tab2 = 23'b00010010000111010100100;
12'd3914 : tab2 = 23'b00010010000000100110100;
12'd3915 : tab2 = 23'b00010001111001111000100;
12'd3916 : tab2 = 23'b00010001110011001011011;
12'd3917 : tab2 = 23'b00010001101100011101101;
12'd3918 : tab2 = 23'b00010001100101110000101;
12'd3919 : tab2 = 23'b00010001011111000011100;
12'd3920 : tab2 = 23'b00010001011000010111010;
12'd3921 : tab2 = 23'b00010001010001101010110;
12'd3922 : tab2 = 23'b00010001001010111110101;
12'd3923 : tab2 = 23'b00010001000100010011000;
12'd3924 : tab2 = 23'b00010000111101100111101;
12'd3925 : tab2 = 23'b00010000110110111100011;
12'd3926 : tab2 = 23'b00010000110000010001100;
12'd3927 : tab2 = 23'b00010000101001100110101;
12'd3928 : tab2 = 23'b00010000100010111100000;
12'd3929 : tab2 = 23'b00010000011100010001111;
12'd3930 : tab2 = 23'b00010000010101101000110;
12'd3931 : tab2 = 23'b00010000001110111110111;
12'd3932 : tab2 = 23'b00010000001000010101011;
12'd3933 : tab2 = 23'b00010000000001101100100;
12'd3934 : tab2 = 23'b00001111111011000011110;
12'd3935 : tab2 = 23'b00001111110100011011011;
12'd3936 : tab2 = 23'b00001111101101110010111;
12'd3937 : tab2 = 23'b00001111100111001011000;
12'd3938 : tab2 = 23'b00001111100000100011100;
12'd3939 : tab2 = 23'b00001111011001111100000;
12'd3940 : tab2 = 23'b00001111010011010100101;
12'd3941 : tab2 = 23'b00001111001100101101111;
12'd3942 : tab2 = 23'b00001111000110000111100;
12'd3943 : tab2 = 23'b00001110111111100000110;
12'd3944 : tab2 = 23'b00001110111000111011000;
12'd3945 : tab2 = 23'b00001110110010010101011;
12'd3946 : tab2 = 23'b00001110101011101111011;
12'd3947 : tab2 = 23'b00001110100101001010010;
12'd3948 : tab2 = 23'b00001110011110100101010;
12'd3949 : tab2 = 23'b00001110011000000000011;
12'd3950 : tab2 = 23'b00001110010001011011110;
12'd3951 : tab2 = 23'b00001110001010110111110;
12'd3952 : tab2 = 23'b00001110000100010100000;
12'd3953 : tab2 = 23'b00001101111101110000100;
12'd3954 : tab2 = 23'b00001101110111001100111;
12'd3955 : tab2 = 23'b00001101110000101001100;
12'd3956 : tab2 = 23'b00001101101010000110111;
12'd3957 : tab2 = 23'b00001101100011100100001;
12'd3958 : tab2 = 23'b00001101011101000010000;
12'd3959 : tab2 = 23'b00001101010110011111111;
12'd3960 : tab2 = 23'b00001101001111111101110;
12'd3961 : tab2 = 23'b00001101001001011100100;
12'd3962 : tab2 = 23'b00001101000010111010111;
12'd3963 : tab2 = 23'b00001100111100011001111;
12'd3964 : tab2 = 23'b00001100110101111001011;
12'd3965 : tab2 = 23'b00001100101111011000101;
12'd3966 : tab2 = 23'b00001100101000111000101;
12'd3967 : tab2 = 23'b00001100100010011000110;
12'd3968 : tab2 = 23'b00001100011011111001000;
12'd3969 : tab2 = 23'b00001100010101011001011;
12'd3970 : tab2 = 23'b00001100001110111001111;
12'd3971 : tab2 = 23'b00001100001000011011001;
12'd3972 : tab2 = 23'b00001100000001111100101;
12'd3973 : tab2 = 23'b00001011111011011110001;
12'd3974 : tab2 = 23'b00001011110100111111110;
12'd3975 : tab2 = 23'b00001011101110100010011;
12'd3976 : tab2 = 23'b00001011101000000100101;
12'd3977 : tab2 = 23'b00001011100001100111000;
12'd3978 : tab2 = 23'b00001011011011001001111;
12'd3979 : tab2 = 23'b00001011010100101100110;
12'd3980 : tab2 = 23'b00001011001110010000101;
12'd3981 : tab2 = 23'b00001011000111110100001;
12'd3982 : tab2 = 23'b00001011000001011000010;
12'd3983 : tab2 = 23'b00001010111010111100010;
12'd3984 : tab2 = 23'b00001010110100100001000;
12'd3985 : tab2 = 23'b00001010101110000101010;
12'd3986 : tab2 = 23'b00001010100111101010100;
12'd3987 : tab2 = 23'b00001010100001001111100;
12'd3988 : tab2 = 23'b00001010011010110101010;
12'd3989 : tab2 = 23'b00001010010100011010110;
12'd3990 : tab2 = 23'b00001010001110000000111;
12'd3991 : tab2 = 23'b00001010000111100110111;
12'd3992 : tab2 = 23'b00001010000001001101100;
12'd3993 : tab2 = 23'b00001001111010110100010;
12'd3994 : tab2 = 23'b00001001110100011011000;
12'd3995 : tab2 = 23'b00001001101110000010101;
12'd3996 : tab2 = 23'b00001001100111101010001;
12'd3997 : tab2 = 23'b00001001100001010001101;
12'd3998 : tab2 = 23'b00001001011010111001101;
12'd3999 : tab2 = 23'b00001001010100100010011;
12'd4000 : tab2 = 23'b00001001001110001010101;
12'd4001 : tab2 = 23'b00001001000111110011011;
12'd4002 : tab2 = 23'b00001001000001011100100;
12'd4003 : tab2 = 23'b00001000111011000110001;
12'd4004 : tab2 = 23'b00001000110100101111100;
12'd4005 : tab2 = 23'b00001000101110011001000;
12'd4006 : tab2 = 23'b00001000101000000011010;
12'd4007 : tab2 = 23'b00001000100001101101110;
12'd4008 : tab2 = 23'b00001000011011011000011;
12'd4009 : tab2 = 23'b00001000010101000011000;
12'd4010 : tab2 = 23'b00001000001110101110000;
12'd4011 : tab2 = 23'b00001000001000011001010;
12'd4012 : tab2 = 23'b00001000000010000101000;
12'd4013 : tab2 = 23'b00000111111011110000110;
12'd4014 : tab2 = 23'b00000111110101011100110;
12'd4015 : tab2 = 23'b00000111101111001001100;
12'd4016 : tab2 = 23'b00000111101000110101101;
12'd4017 : tab2 = 23'b00000111100010100010101;
12'd4018 : tab2 = 23'b00000111011100001111110;
12'd4019 : tab2 = 23'b00000111010101111100110;
12'd4020 : tab2 = 23'b00000111001111101010111;
12'd4021 : tab2 = 23'b00000111001001011000101;
12'd4022 : tab2 = 23'b00000111000011000110111;
12'd4023 : tab2 = 23'b00000110111100110100111;
12'd4024 : tab2 = 23'b00000110110110100011101;
12'd4025 : tab2 = 23'b00000110110000010010101;
12'd4026 : tab2 = 23'b00000110101010000001100;
12'd4027 : tab2 = 23'b00000110100011110000110;
12'd4028 : tab2 = 23'b00000110011101100000011;
12'd4029 : tab2 = 23'b00000110010111010000001;
12'd4030 : tab2 = 23'b00000110010001000000100;
12'd4031 : tab2 = 23'b00000110001010110000111;
12'd4032 : tab2 = 23'b00000110000100100001010;
12'd4033 : tab2 = 23'b00000101111110010010001;
12'd4034 : tab2 = 23'b00000101111000000011001;
12'd4035 : tab2 = 23'b00000101110001110100111;
12'd4036 : tab2 = 23'b00000101101011100110000;
12'd4037 : tab2 = 23'b00000101100101011000000;
12'd4038 : tab2 = 23'b00000101011111001010001;
12'd4039 : tab2 = 23'b00000101011000111100011;
12'd4040 : tab2 = 23'b00000101010010101110110;
12'd4041 : tab2 = 23'b00000101001100100001111;
12'd4042 : tab2 = 23'b00000101000110010100110;
12'd4043 : tab2 = 23'b00000101000000000111110;
12'd4044 : tab2 = 23'b00000100111001111011010;
12'd4045 : tab2 = 23'b00000100110011101111101;
12'd4046 : tab2 = 23'b00000100101101100011010;
12'd4047 : tab2 = 23'b00000100100111010111101;
12'd4048 : tab2 = 23'b00000100100001001100000;
12'd4049 : tab2 = 23'b00000100011011000001000;
12'd4050 : tab2 = 23'b00000100010100110101111;
12'd4051 : tab2 = 23'b00000100001110101011010;
12'd4052 : tab2 = 23'b00000100001000100000100;
12'd4053 : tab2 = 23'b00000100000010010110011;
12'd4054 : tab2 = 23'b00000011111100001100011;
12'd4055 : tab2 = 23'b00000011110110000010011;
12'd4056 : tab2 = 23'b00000011101111111001000;
12'd4057 : tab2 = 23'b00000011101001101111101;
12'd4058 : tab2 = 23'b00000011100011100110101;
12'd4059 : tab2 = 23'b00000011011101011101111;
12'd4060 : tab2 = 23'b00000011010111010101010;
12'd4061 : tab2 = 23'b00000011010001001101000;
12'd4062 : tab2 = 23'b00000011001011000100111;
12'd4063 : tab2 = 23'b00000011000100111101010;
12'd4064 : tab2 = 23'b00000010111110110101100;
12'd4065 : tab2 = 23'b00000010111000101110010;
12'd4066 : tab2 = 23'b00000010110010100110110;
12'd4067 : tab2 = 23'b00000010101100100000000;
12'd4068 : tab2 = 23'b00000010100110011001011;
12'd4069 : tab2 = 23'b00000010100000010010111;
12'd4070 : tab2 = 23'b00000010011010001100111;
12'd4071 : tab2 = 23'b00000010010100000111010;
12'd4072 : tab2 = 23'b00000010001110000001001;
12'd4073 : tab2 = 23'b00000010000111111011101;
12'd4074 : tab2 = 23'b00000010000001110110100;
12'd4075 : tab2 = 23'b00000001111011110001111;
12'd4076 : tab2 = 23'b00000001110101101101000;
12'd4077 : tab2 = 23'b00000001101111101000001;
12'd4078 : tab2 = 23'b00000001101001100100010;
12'd4079 : tab2 = 23'b00000001100011100000011;
12'd4080 : tab2 = 23'b00000001011101011100100;
12'd4081 : tab2 = 23'b00000001010111011000111;
12'd4082 : tab2 = 23'b00000001010001010101011;
12'd4083 : tab2 = 23'b00000001001011010010101;
12'd4084 : tab2 = 23'b00000001000101001111101;
12'd4085 : tab2 = 23'b00000000111111001101001;
12'd4086 : tab2 = 23'b00000000111001001011000;
12'd4087 : tab2 = 23'b00000000110011001000101;
12'd4088 : tab2 = 23'b00000000101101000110110;
12'd4089 : tab2 = 23'b00000000100111000101000;
12'd4090 : tab2 = 23'b00000000100001000011110;
12'd4091 : tab2 = 23'b00000000011011000010100;
12'd4092 : tab2 = 23'b00000000010101000001011;
12'd4093 : tab2 = 23'b00000000001111000001001;
12'd4094 : tab2 = 23'b00000000001001000000100;
12'd4095 : tab2 = 23'b00000000000011000000000;
  endcase
  end
  endfunction


  wire [0:0] swire5;
  wire [7:0] ewire5;
  wire [22:0] mwire5;

  assign swire5 = x[31];
  assign ewire5 = x[30:23];
  assign mwire5 = x[22:0];

  wire [23:0] mawire5;
  wire [7:0] eawire5;

  assign mawire5 = (ewire5 == 8'b0) ? {1'b0,mwire5[22:0]} : {1'b1,mwire5[22:0]};
  assign eawire5 = ((ewire5+1) >> 1) + 8'd63 + (&{~ewire5[0],mwire5});


  reg [0:0] swirereg4;
  reg [7:0] ewirereg4;
  reg [22:0] mwirereg4;
  reg [23:0] mawirereg4;
  reg [7:0] eawirereg4;
  reg [0:0] swirereg3;
  reg [7:0] ewirereg3;
  reg [22:0] mwirereg3;
  reg [23:0] mawirereg3;
  reg [7:0] eawirereg3;


  wire [23:0] nibunno3xwire5;
  reg [23:0] nibunno3xreg4;
  reg [23:0] nibunno3xreg3;
  
  assign nibunno3xwire5 = {1'b1,tab({~ewire5[0],mwire5[22:12]})};

  wire [23:0] nibunnox3wire5;
  reg [23:0] nibunnox3reg4;
  
  assign nibunnox3wire5 = {1'b1,tab2({~ewire5[0],mwire5[22:12]})};

  wire [47:0] nibunnox3awire4;
  reg [47:0] nibunnox3areg3;
  //////////
  assign nibunnox3awire4 = mawirereg4 * nibunnox3reg4;
////////
  wire [47:0] nibunnox3ak1;
  wire [47:0] nibunnox3ak0;
  assign nibunnox3ak1 = (ewirereg3[0] == 1) ? (({~ewirereg3[0],mwirereg3[22:12]} > 12'd1202) ? (nibunnox3areg3 >> 2) : nibunnox3areg3 >> 1) : ( ({~ewirereg3[0],mwirereg3[22:12]} > 12'd2579) ? (nibunnox3areg3 >> 2) : (nibunnox3areg3 >> 1));
  assign nibunnox3ak0 = ({~ewirereg3[0],mwirereg3[22:12]} > 12'd2303) ? (nibunnox3ak1 << 1) : nibunnox3ak1;
  
  wire [23:0] nibunnox3ak;
  wire [23:0] rootabunno1wire3;
  wire [47:0] rootawire2;

  reg [23:0] rootabunno1reg2;
  reg [47:0] rootareg;

  reg [0:0] swirereg2;
  reg [7:0] ewirereg2;
  reg [23:0] mawirereg2;
  reg [7:0] eawirereg2;

  assign nibunnox3ak = {nibunnox3ak0[47:24]};
  assign rootabunno1wire3 = nibunno3xreg3 - nibunnox3ak;
///////
  assign rootawire2 = mawirereg2 * rootabunno1reg2;

  reg [0:0] swirereg;
  reg [7:0] ewirereg;
  reg [7:0] eawirereg;
////

  wire [47:0] keta;
  wire [22:0] ans;
  
  assign keta = (rootareg[47] == 0) ?
               ((rootareg[46] == 0) ?
               ((rootareg[45] == 0) ? 
               ((rootareg[44] == 0) ? (rootareg << 5) : (rootareg << 4)) : (rootareg << 3)) : (rootareg << 2)): (rootareg << 1);
  assign ans = keta[47:25];
  assign y = (ewirereg == 23'b0 || ewirereg == 23'd255) ? {swirereg,31'b0} : {swirereg,eawirereg,ans} ;

  always @(posedge clk) begin
    
    swirereg4<=swire5;
    ewirereg4<=ewire5;
    mwirereg4<=mwire5;
    mawirereg4<=mawire5;
    eawirereg4<=eawire5;
    swirereg3<=swirereg4;
    ewirereg3<=ewirereg4;
    mwirereg3<=mwirereg4;
    mawirereg3<=mawirereg4;
    eawirereg3<=eawirereg4;
    nibunno3xreg4<=nibunno3xwire5;
    nibunno3xreg3<=nibunno3xreg4;
    nibunnox3reg4<=nibunnox3wire5;
    nibunnox3areg3<=nibunnox3awire4;
    rootabunno1reg2<=rootabunno1wire3;
    rootareg<=rootawire2;
    swirereg2<=swirereg3;
    ewirereg2<=ewirereg3;
    mawirereg2<=mawirereg3;
    eawirereg2<=eawirereg3;
    swirereg<=swirereg2;
    ewirereg<=ewirereg2;
    eawirereg<=eawirereg2;
  end
  
endmodule
`default_nettype wire

