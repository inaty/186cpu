`timescale 1ns / 1ps
`default_nettype none

module finv_d(
  input wire [31:0] x,
  output wire [31:0] y,
  input wire clk);

  function [22:0] tab (
    input [10:0] M
  );
  begin
  case(M)
11'd0 : tab = 23'b11111111111000000000011;
11'd1 : tab = 23'b11111111101000000001011;
11'd2 : tab = 23'b11111111011000000011011;
11'd3 : tab = 23'b11111111001000000110011;
11'd4 : tab = 23'b11111110111000001010011;
11'd5 : tab = 23'b11111110101000001111011;
11'd6 : tab = 23'b11111110011000010101010;
11'd7 : tab = 23'b11111110001000011100010;
11'd8 : tab = 23'b11111101111000100100010;
11'd9 : tab = 23'b11111101101000101101010;
11'd10 : tab = 23'b11111101011000110111000;
11'd11 : tab = 23'b11111101001001000010000;
11'd12 : tab = 23'b11111100111001001110000;
11'd13 : tab = 23'b11111100101001011010110;
11'd14 : tab = 23'b11111100011001101000101;
11'd15 : tab = 23'b11111100001001110111100;
11'd16 : tab = 23'b11111011111010000111010;
11'd17 : tab = 23'b11111011101010011000000;
11'd18 : tab = 23'b11111011011010101001111;
11'd19 : tab = 23'b11111011001010111100100;
11'd20 : tab = 23'b11111010111011010000010;
11'd21 : tab = 23'b11111010101011100101000;
11'd22 : tab = 23'b11111010011011111010100;
11'd23 : tab = 23'b11111010001100010001010;
11'd24 : tab = 23'b11111001111100101000110;
11'd25 : tab = 23'b11111001101101000001011;
11'd26 : tab = 23'b11111001011101011010111;
11'd27 : tab = 23'b11111001001101110101011;
11'd28 : tab = 23'b11111000111110010000110;
11'd29 : tab = 23'b11111000101110101101010;
11'd30 : tab = 23'b11111000011111001010100;
11'd31 : tab = 23'b11111000001111101000111;
11'd32 : tab = 23'b11111000000000001000001;
11'd33 : tab = 23'b11110111110000101000010;
11'd34 : tab = 23'b11110111100001001001100;
11'd35 : tab = 23'b11110111010001101011101;
11'd36 : tab = 23'b11110111000010001110110;
11'd37 : tab = 23'b11110110110010110010110;
11'd38 : tab = 23'b11110110100011010111110;
11'd39 : tab = 23'b11110110010011111101100;
11'd40 : tab = 23'b11110110000100100100100;
11'd41 : tab = 23'b11110101110101001100010;
11'd42 : tab = 23'b11110101100101110101000;
11'd43 : tab = 23'b11110101010110011110110;
11'd44 : tab = 23'b11110101000111001001010;
11'd45 : tab = 23'b11110100110111110100111;
11'd46 : tab = 23'b11110100101000100001011;
11'd47 : tab = 23'b11110100011001001110110;
11'd48 : tab = 23'b11110100001001111101001;
11'd49 : tab = 23'b11110011111010101100100;
11'd50 : tab = 23'b11110011101011011100110;
11'd51 : tab = 23'b11110011011100001101110;
11'd52 : tab = 23'b11110011001100111111111;
11'd53 : tab = 23'b11110010111101110011000;
11'd54 : tab = 23'b11110010101110100110110;
11'd55 : tab = 23'b11110010011111011011110;
11'd56 : tab = 23'b11110010010000010001100;
11'd57 : tab = 23'b11110010000001001000010;
11'd58 : tab = 23'b11110001110001111111110;
11'd59 : tab = 23'b11110001100010111000011;
11'd60 : tab = 23'b11110001010011110001110;
11'd61 : tab = 23'b11110001000100101100010;
11'd62 : tab = 23'b11110000110101100111100;
11'd63 : tab = 23'b11110000100110100011110;
11'd64 : tab = 23'b11110000010111100000111;
11'd65 : tab = 23'b11110000001000011110111;
11'd66 : tab = 23'b11101111111001011101110;
11'd67 : tab = 23'b11101111101010011101101;
11'd68 : tab = 23'b11101111011011011110100;
11'd69 : tab = 23'b11101111001100100000000;
11'd70 : tab = 23'b11101110111101100010101;
11'd71 : tab = 23'b11101110101110100110001;
11'd72 : tab = 23'b11101110011111101010100;
11'd73 : tab = 23'b11101110010000101111110;
11'd74 : tab = 23'b11101110000001110110000;
11'd75 : tab = 23'b11101101110010111101000;
11'd76 : tab = 23'b11101101100100000101000;
11'd77 : tab = 23'b11101101010101001101111;
11'd78 : tab = 23'b11101101000110010111101;
11'd79 : tab = 23'b11101100110111100010010;
11'd80 : tab = 23'b11101100101000101101110;
11'd81 : tab = 23'b11101100011001111010010;
11'd82 : tab = 23'b11101100001011000111101;
11'd83 : tab = 23'b11101011111100010101110;
11'd84 : tab = 23'b11101011101101100100111;
11'd85 : tab = 23'b11101011011110110100111;
11'd86 : tab = 23'b11101011010000000101110;
11'd87 : tab = 23'b11101011000001010111100;
11'd88 : tab = 23'b11101010110010101010001;
11'd89 : tab = 23'b11101010100011111101101;
11'd90 : tab = 23'b11101010010101010010000;
11'd91 : tab = 23'b11101010000110100111010;
11'd92 : tab = 23'b11101001110111111101100;
11'd93 : tab = 23'b11101001101001010100100;
11'd94 : tab = 23'b11101001011010101100011;
11'd95 : tab = 23'b11101001001100000101010;
11'd96 : tab = 23'b11101000111101011110110;
11'd97 : tab = 23'b11101000101110111001011;
11'd98 : tab = 23'b11101000100000010100110;
11'd99 : tab = 23'b11101000010001110001000;
11'd100 : tab = 23'b11101000000011001110001;
11'd101 : tab = 23'b11100111110100101100000;
11'd102 : tab = 23'b11100111100110001011000;
11'd103 : tab = 23'b11100111010111101010110;
11'd104 : tab = 23'b11100111001001001011010;
11'd105 : tab = 23'b11100110111010101100110;
11'd106 : tab = 23'b11100110101100001111000;
11'd107 : tab = 23'b11100110011101110010010;
11'd108 : tab = 23'b11100110001111010110010;
11'd109 : tab = 23'b11100110000000111011000;
11'd110 : tab = 23'b11100101110010100000110;
11'd111 : tab = 23'b11100101100100000111011;
11'd112 : tab = 23'b11100101010101101110110;
11'd113 : tab = 23'b11100101000111010111001;
11'd114 : tab = 23'b11100100111001000000010;
11'd115 : tab = 23'b11100100101010101010010;
11'd116 : tab = 23'b11100100011100010101001;
11'd117 : tab = 23'b11100100001110000000110;
11'd118 : tab = 23'b11100011111111101101010;
11'd119 : tab = 23'b11100011110001011010110;
11'd120 : tab = 23'b11100011100011001001000;
11'd121 : tab = 23'b11100011010100111000000;
11'd122 : tab = 23'b11100011000110100111111;
11'd123 : tab = 23'b11100010111000011000101;
11'd124 : tab = 23'b11100010101010001010010;
11'd125 : tab = 23'b11100010011011111100101;
11'd126 : tab = 23'b11100010001101101111111;
11'd127 : tab = 23'b11100001111111100100000;
11'd128 : tab = 23'b11100001110001011000111;
11'd129 : tab = 23'b11100001100011001110110;
11'd130 : tab = 23'b11100001010101000101010;
11'd131 : tab = 23'b11100001000110111100110;
11'd132 : tab = 23'b11100000111000110101000;
11'd133 : tab = 23'b11100000101010101110000;
11'd134 : tab = 23'b11100000011100101000000;
11'd135 : tab = 23'b11100000001110100010110;
11'd136 : tab = 23'b11100000000000011110010;
11'd137 : tab = 23'b11011111110010011010101;
11'd138 : tab = 23'b11011111100100010111110;
11'd139 : tab = 23'b11011111010110010101110;
11'd140 : tab = 23'b11011111001000010100110;
11'd141 : tab = 23'b11011110111010010100011;
11'd142 : tab = 23'b11011110101100010100110;
11'd143 : tab = 23'b11011110011110010110001;
11'd144 : tab = 23'b11011110010000011000010;
11'd145 : tab = 23'b11011110000010011011010;
11'd146 : tab = 23'b11011101110100011111000;
11'd147 : tab = 23'b11011101100110100011100;
11'd148 : tab = 23'b11011101011000101000111;
11'd149 : tab = 23'b11011101001010101111000;
11'd150 : tab = 23'b11011100111100110110000;
11'd151 : tab = 23'b11011100101110111101111;
11'd152 : tab = 23'b11011100100001000110100;
11'd153 : tab = 23'b11011100010011001111111;
11'd154 : tab = 23'b11011100000101011010001;
11'd155 : tab = 23'b11011011110111100101010;
11'd156 : tab = 23'b11011011101001110001000;
11'd157 : tab = 23'b11011011011011111101101;
11'd158 : tab = 23'b11011011001110001011000;
11'd159 : tab = 23'b11011011000000011001010;
11'd160 : tab = 23'b11011010110010101000010;
11'd161 : tab = 23'b11011010100100111000001;
11'd162 : tab = 23'b11011010010111001000110;
11'd163 : tab = 23'b11011010001001011010001;
11'd164 : tab = 23'b11011001111011101100011;
11'd165 : tab = 23'b11011001101101111111010;
11'd166 : tab = 23'b11011001100000010011010;
11'd167 : tab = 23'b11011001010010100111110;
11'd168 : tab = 23'b11011001000100111101001;
11'd169 : tab = 23'b11011000110111010011010;
11'd170 : tab = 23'b11011000101001101010010;
11'd171 : tab = 23'b11011000011100000010000;
11'd172 : tab = 23'b11011000001110011010100;
11'd173 : tab = 23'b11011000000000110011110;
11'd174 : tab = 23'b11010111110011001110000;
11'd175 : tab = 23'b11010111100101101000110;
11'd176 : tab = 23'b11010111011000000100100;
11'd177 : tab = 23'b11010111001010100000111;
11'd178 : tab = 23'b11010110111100111110001;
11'd179 : tab = 23'b11010110101111011100001;
11'd180 : tab = 23'b11010110100001111011000;
11'd181 : tab = 23'b11010110010100011010100;
11'd182 : tab = 23'b11010110000110111010110;
11'd183 : tab = 23'b11010101111001011011111;
11'd184 : tab = 23'b11010101101011111101110;
11'd185 : tab = 23'b11010101011110100000011;
11'd186 : tab = 23'b11010101010001000011110;
11'd187 : tab = 23'b11010101000011101000000;
11'd188 : tab = 23'b11010100110110001101000;
11'd189 : tab = 23'b11010100101000110010110;
11'd190 : tab = 23'b11010100011011011001001;
11'd191 : tab = 23'b11010100001110000000100;
11'd192 : tab = 23'b11010100000000101000100;
11'd193 : tab = 23'b11010011110011010001010;
11'd194 : tab = 23'b11010011100101111010110;
11'd195 : tab = 23'b11010011011000100101000;
11'd196 : tab = 23'b11010011001011010000001;
11'd197 : tab = 23'b11010010111101111100000;
11'd198 : tab = 23'b11010010110000101000100;
11'd199 : tab = 23'b11010010100011010101111;
11'd200 : tab = 23'b11010010010110000100000;
11'd201 : tab = 23'b11010010001000110010110;
11'd202 : tab = 23'b11010001111011100010100;
11'd203 : tab = 23'b11010001101110010010110;
11'd204 : tab = 23'b11010001100001000100000;
11'd205 : tab = 23'b11010001010011110101110;
11'd206 : tab = 23'b11010001000110101000100;
11'd207 : tab = 23'b11010000111001011011110;
11'd208 : tab = 23'b11010000101100001111111;
11'd209 : tab = 23'b11010000011111000100110;
11'd210 : tab = 23'b11010000010001111010011;
11'd211 : tab = 23'b11010000000100110000110;
11'd212 : tab = 23'b11001111110111100111110;
11'd213 : tab = 23'b11001111101010011111110;
11'd214 : tab = 23'b11001111011101011000010;
11'd215 : tab = 23'b11001111010000010001101;
11'd216 : tab = 23'b11001111000011001011110;
11'd217 : tab = 23'b11001110110110000110100;
11'd218 : tab = 23'b11001110101001000010000;
11'd219 : tab = 23'b11001110011011111110010;
11'd220 : tab = 23'b11001110001110111011010;
11'd221 : tab = 23'b11001110000001111001001;
11'd222 : tab = 23'b11001101110100110111101;
11'd223 : tab = 23'b11001101100111110110111;
11'd224 : tab = 23'b11001101011010110110110;
11'd225 : tab = 23'b11001101001101110111100;
11'd226 : tab = 23'b11001101000000111000111;
11'd227 : tab = 23'b11001100110011111011000;
11'd228 : tab = 23'b11001100100110111110000;
11'd229 : tab = 23'b11001100011010000001100;
11'd230 : tab = 23'b11001100001101000110000;
11'd231 : tab = 23'b11001100000000001011000;
11'd232 : tab = 23'b11001011110011010000110;
11'd233 : tab = 23'b11001011100110010111010;
11'd234 : tab = 23'b11001011011001011110100;
11'd235 : tab = 23'b11001011001100100110100;
11'd236 : tab = 23'b11001010111111101111001;
11'd237 : tab = 23'b11001010110010111000100;
11'd238 : tab = 23'b11001010100110000010110;
11'd239 : tab = 23'b11001010011001001101100;
11'd240 : tab = 23'b11001010001100011001000;
11'd241 : tab = 23'b11001001111111100101011;
11'd242 : tab = 23'b11001001110010110010011;
11'd243 : tab = 23'b11001001100110000000000;
11'd244 : tab = 23'b11001001011001001110100;
11'd245 : tab = 23'b11001001001100011101101;
11'd246 : tab = 23'b11001000111111101101100;
11'd247 : tab = 23'b11001000110010111110000;
11'd248 : tab = 23'b11001000100110001111010;
11'd249 : tab = 23'b11001000011001100001010;
11'd250 : tab = 23'b11001000001100110011111;
11'd251 : tab = 23'b11001000000000000111010;
11'd252 : tab = 23'b11000111110011011011100;
11'd253 : tab = 23'b11000111100110110000010;
11'd254 : tab = 23'b11000111011010000101110;
11'd255 : tab = 23'b11000111001101011011111;
11'd256 : tab = 23'b11000111000000110010111;
11'd257 : tab = 23'b11000110110100001010100;
11'd258 : tab = 23'b11000110100111100010110;
11'd259 : tab = 23'b11000110011010111011110;
11'd260 : tab = 23'b11000110001110010101100;
11'd261 : tab = 23'b11000110000001110000000;
11'd262 : tab = 23'b11000101110101001011000;
11'd263 : tab = 23'b11000101101000100110110;
11'd264 : tab = 23'b11000101011100000011011;
11'd265 : tab = 23'b11000101001111100000100;
11'd266 : tab = 23'b11000101000010111110100;
11'd267 : tab = 23'b11000100110110011101000;
11'd268 : tab = 23'b11000100101001111100010;
11'd269 : tab = 23'b11000100011101011100010;
11'd270 : tab = 23'b11000100010000111101000;
11'd271 : tab = 23'b11000100000100011110010;
11'd272 : tab = 23'b11000011111000000000010;
11'd273 : tab = 23'b11000011101011100011000;
11'd274 : tab = 23'b11000011011111000110100;
11'd275 : tab = 23'b11000011010010101010100;
11'd276 : tab = 23'b11000011000110001111010;
11'd277 : tab = 23'b11000010111001110100110;
11'd278 : tab = 23'b11000010101101011011000;
11'd279 : tab = 23'b11000010100001000001110;
11'd280 : tab = 23'b11000010010100101001010;
11'd281 : tab = 23'b11000010001000010001100;
11'd282 : tab = 23'b11000001111011111010010;
11'd283 : tab = 23'b11000001101111100011111;
11'd284 : tab = 23'b11000001100011001110001;
11'd285 : tab = 23'b11000001010110111001000;
11'd286 : tab = 23'b11000001001010100100100;
11'd287 : tab = 23'b11000000111110010000110;
11'd288 : tab = 23'b11000000110001111101110;
11'd289 : tab = 23'b11000000100101101011010;
11'd290 : tab = 23'b11000000011001011001101;
11'd291 : tab = 23'b11000000001101001000100;
11'd292 : tab = 23'b11000000000000111000010;
11'd293 : tab = 23'b10111111110100101000100;
11'd294 : tab = 23'b10111111101000011001011;
11'd295 : tab = 23'b10111111011100001011000;
11'd296 : tab = 23'b10111111001111111101010;
11'd297 : tab = 23'b10111111000011110000010;
11'd298 : tab = 23'b10111110110111100100000;
11'd299 : tab = 23'b10111110101011011000010;
11'd300 : tab = 23'b10111110011111001101001;
11'd301 : tab = 23'b10111110010011000010110;
11'd302 : tab = 23'b10111110000110111001000;
11'd303 : tab = 23'b10111101111010110000000;
11'd304 : tab = 23'b10111101101110100111100;
11'd305 : tab = 23'b10111101100010011111111;
11'd306 : tab = 23'b10111101010110011000110;
11'd307 : tab = 23'b10111101001010010010010;
11'd308 : tab = 23'b10111100111110001100101;
11'd309 : tab = 23'b10111100110010000111100;
11'd310 : tab = 23'b10111100100110000011000;
11'd311 : tab = 23'b10111100011001111111010;
11'd312 : tab = 23'b10111100001101111100000;
11'd313 : tab = 23'b10111100000001111001101;
11'd314 : tab = 23'b10111011110101110111110;
11'd315 : tab = 23'b10111011101001110110100;
11'd316 : tab = 23'b10111011011101110110000;
11'd317 : tab = 23'b10111011010001110110010;
11'd318 : tab = 23'b10111011000101110110111;
11'd319 : tab = 23'b10111010111001111000010;
11'd320 : tab = 23'b10111010101101111010011;
11'd321 : tab = 23'b10111010100001111101000;
11'd322 : tab = 23'b10111010010110000000100;
11'd323 : tab = 23'b10111010001010000100011;
11'd324 : tab = 23'b10111001111110001001000;
11'd325 : tab = 23'b10111001110010001110010;
11'd326 : tab = 23'b10111001100110010100010;
11'd327 : tab = 23'b10111001011010011010110;
11'd328 : tab = 23'b10111001001110100010000;
11'd329 : tab = 23'b10111001000010101001111;
11'd330 : tab = 23'b10111000110110110010011;
11'd331 : tab = 23'b10111000101010111011100;
11'd332 : tab = 23'b10111000011111000101010;
11'd333 : tab = 23'b10111000010011001111101;
11'd334 : tab = 23'b10111000000111011010110;
11'd335 : tab = 23'b10110111111011100110010;
11'd336 : tab = 23'b10110111101111110010101;
11'd337 : tab = 23'b10110111100011111111100;
11'd338 : tab = 23'b10110111011000001101001;
11'd339 : tab = 23'b10110111001100011011011;
11'd340 : tab = 23'b10110111000000101010010;
11'd341 : tab = 23'b10110110110100111001101;
11'd342 : tab = 23'b10110110101001001001110;
11'd343 : tab = 23'b10110110011101011010100;
11'd344 : tab = 23'b10110110010001101011110;
11'd345 : tab = 23'b10110110000101111101110;
11'd346 : tab = 23'b10110101111010010000100;
11'd347 : tab = 23'b10110101101110100011101;
11'd348 : tab = 23'b10110101100010110111100;
11'd349 : tab = 23'b10110101010111001100000;
11'd350 : tab = 23'b10110101001011100001000;
11'd351 : tab = 23'b10110100111111110110110;
11'd352 : tab = 23'b10110100110100001101001;
11'd353 : tab = 23'b10110100101000100100001;
11'd354 : tab = 23'b10110100011100111011110;
11'd355 : tab = 23'b10110100010001010011111;
11'd356 : tab = 23'b10110100000101101100110;
11'd357 : tab = 23'b10110011111010000110010;
11'd358 : tab = 23'b10110011101110100000010;
11'd359 : tab = 23'b10110011100010111010111;
11'd360 : tab = 23'b10110011010111010110010;
11'd361 : tab = 23'b10110011001011110010000;
11'd362 : tab = 23'b10110011000000001110101;
11'd363 : tab = 23'b10110010110100101011110;
11'd364 : tab = 23'b10110010101001001001100;
11'd365 : tab = 23'b10110010011101100111110;
11'd366 : tab = 23'b10110010010010000110110;
11'd367 : tab = 23'b10110010000110100110011;
11'd368 : tab = 23'b10110001111011000110100;
11'd369 : tab = 23'b10110001101111100111011;
11'd370 : tab = 23'b10110001100100001000110;
11'd371 : tab = 23'b10110001011000101010110;
11'd372 : tab = 23'b10110001001101001101100;
11'd373 : tab = 23'b10110001000001110000101;
11'd374 : tab = 23'b10110000110110010100100;
11'd375 : tab = 23'b10110000101010111001000;
11'd376 : tab = 23'b10110000011111011110000;
11'd377 : tab = 23'b10110000010100000011100;
11'd378 : tab = 23'b10110000001000101001111;
11'd379 : tab = 23'b10101111111101010000110;
11'd380 : tab = 23'b10101111110001111000001;
11'd381 : tab = 23'b10101111100110100000001;
11'd382 : tab = 23'b10101111011011001000110;
11'd383 : tab = 23'b10101111001111110010000;
11'd384 : tab = 23'b10101111000100011011111;
11'd385 : tab = 23'b10101110111001000110010;
11'd386 : tab = 23'b10101110101101110001011;
11'd387 : tab = 23'b10101110100010011101000;
11'd388 : tab = 23'b10101110010111001001010;
11'd389 : tab = 23'b10101110001011110110000;
11'd390 : tab = 23'b10101110000000100011100;
11'd391 : tab = 23'b10101101110101010001100;
11'd392 : tab = 23'b10101101101010000000000;
11'd393 : tab = 23'b10101101011110101111010;
11'd394 : tab = 23'b10101101010011011111000;
11'd395 : tab = 23'b10101101001000001111010;
11'd396 : tab = 23'b10101100111101000000010;
11'd397 : tab = 23'b10101100110001110001111;
11'd398 : tab = 23'b10101100100110100100000;
11'd399 : tab = 23'b10101100011011010110110;
11'd400 : tab = 23'b10101100010000001010000;
11'd401 : tab = 23'b10101100000100111101111;
11'd402 : tab = 23'b10101011111001110010011;
11'd403 : tab = 23'b10101011101110100111011;
11'd404 : tab = 23'b10101011100011011101000;
11'd405 : tab = 23'b10101011011000010011010;
11'd406 : tab = 23'b10101011001101001010000;
11'd407 : tab = 23'b10101011000010000001100;
11'd408 : tab = 23'b10101010110110111001011;
11'd409 : tab = 23'b10101010101011110010000;
11'd410 : tab = 23'b10101010100000101011000;
11'd411 : tab = 23'b10101010010101100100110;
11'd412 : tab = 23'b10101010001010011111000;
11'd413 : tab = 23'b10101001111111011001111;
11'd414 : tab = 23'b10101001110100010101010;
11'd415 : tab = 23'b10101001101001010001010;
11'd416 : tab = 23'b10101001011110001101111;
11'd417 : tab = 23'b10101001010011001011000;
11'd418 : tab = 23'b10101001001000001000110;
11'd419 : tab = 23'b10101000111101000111001;
11'd420 : tab = 23'b10101000110010000110000;
11'd421 : tab = 23'b10101000100111000101011;
11'd422 : tab = 23'b10101000011100000101011;
11'd423 : tab = 23'b10101000010001000110000;
11'd424 : tab = 23'b10101000000110000111001;
11'd425 : tab = 23'b10100111111011001000110;
11'd426 : tab = 23'b10100111110000001011001;
11'd427 : tab = 23'b10100111100101001110000;
11'd428 : tab = 23'b10100111011010010001100;
11'd429 : tab = 23'b10100111001111010101011;
11'd430 : tab = 23'b10100111000100011001111;
11'd431 : tab = 23'b10100110111001011111000;
11'd432 : tab = 23'b10100110101110100100110;
11'd433 : tab = 23'b10100110100011101011000;
11'd434 : tab = 23'b10100110011000110001110;
11'd435 : tab = 23'b10100110001101111001001;
11'd436 : tab = 23'b10100110000011000001000;
11'd437 : tab = 23'b10100101111000001001100;
11'd438 : tab = 23'b10100101101101010010101;
11'd439 : tab = 23'b10100101100010011100010;
11'd440 : tab = 23'b10100101010111100110010;
11'd441 : tab = 23'b10100101001100110001000;
11'd442 : tab = 23'b10100101000001111100010;
11'd443 : tab = 23'b10100100110111001000001;
11'd444 : tab = 23'b10100100101100010100100;
11'd445 : tab = 23'b10100100100001100001100;
11'd446 : tab = 23'b10100100010110101111000;
11'd447 : tab = 23'b10100100001011111101000;
11'd448 : tab = 23'b10100100000001001011101;
11'd449 : tab = 23'b10100011110110011010110;
11'd450 : tab = 23'b10100011101011101010100;
11'd451 : tab = 23'b10100011100000111010110;
11'd452 : tab = 23'b10100011010110001011100;
11'd453 : tab = 23'b10100011001011011100111;
11'd454 : tab = 23'b10100011000000101110110;
11'd455 : tab = 23'b10100010110110000001010;
11'd456 : tab = 23'b10100010101011010100010;
11'd457 : tab = 23'b10100010100000100111110;
11'd458 : tab = 23'b10100010010101111011111;
11'd459 : tab = 23'b10100010001011010000100;
11'd460 : tab = 23'b10100010000000100101110;
11'd461 : tab = 23'b10100001110101111011100;
11'd462 : tab = 23'b10100001101011010001110;
11'd463 : tab = 23'b10100001100000101000100;
11'd464 : tab = 23'b10100001010101111111111;
11'd465 : tab = 23'b10100001001011010111110;
11'd466 : tab = 23'b10100001000000110000010;
11'd467 : tab = 23'b10100000110110001001010;
11'd468 : tab = 23'b10100000101011100010110;
11'd469 : tab = 23'b10100000100000111100110;
11'd470 : tab = 23'b10100000010110010111011;
11'd471 : tab = 23'b10100000001011110010100;
11'd472 : tab = 23'b10100000000001001110010;
11'd473 : tab = 23'b10011111110110101010010;
11'd474 : tab = 23'b10011111101100000111001;
11'd475 : tab = 23'b10011111100001100100011;
11'd476 : tab = 23'b10011111010111000010010;
11'd477 : tab = 23'b10011111001100100000100;
11'd478 : tab = 23'b10011111000001111111100;
11'd479 : tab = 23'b10011110110111011110110;
11'd480 : tab = 23'b10011110101100111110110;
11'd481 : tab = 23'b10011110100010011111010;
11'd482 : tab = 23'b10011110011000000000010;
11'd483 : tab = 23'b10011110001101100001110;
11'd484 : tab = 23'b10011110000011000011111;
11'd485 : tab = 23'b10011101111000100110100;
11'd486 : tab = 23'b10011101101110001001100;
11'd487 : tab = 23'b10011101100011101101010;
11'd488 : tab = 23'b10011101011001010001100;
11'd489 : tab = 23'b10011101001110110110000;
11'd490 : tab = 23'b10011101000100011011010;
11'd491 : tab = 23'b10011100111010000001000;
11'd492 : tab = 23'b10011100101111100111011;
11'd493 : tab = 23'b10011100100101001110001;
11'd494 : tab = 23'b10011100011010110101100;
11'd495 : tab = 23'b10011100010000011101011;
11'd496 : tab = 23'b10011100000110000101110;
11'd497 : tab = 23'b10011011111011101110101;
11'd498 : tab = 23'b10011011110001011000000;
11'd499 : tab = 23'b10011011100111000010000;
11'd500 : tab = 23'b10011011011100101100100;
11'd501 : tab = 23'b10011011010010010111010;
11'd502 : tab = 23'b10011011001000000010110;
11'd503 : tab = 23'b10011010111101101110111;
11'd504 : tab = 23'b10011010110011011011011;
11'd505 : tab = 23'b10011010101001001000100;
11'd506 : tab = 23'b10011010011110110110000;
11'd507 : tab = 23'b10011010010100100100000;
11'd508 : tab = 23'b10011010001010010010101;
11'd509 : tab = 23'b10011010000000000001110;
11'd510 : tab = 23'b10011001110101110001011;
11'd511 : tab = 23'b10011001101011100001100;
11'd512 : tab = 23'b10011001100001010010001;
11'd513 : tab = 23'b10011001010111000011010;
11'd514 : tab = 23'b10011001001100110101000;
11'd515 : tab = 23'b10011001000010100111001;
11'd516 : tab = 23'b10011000111000011001110;
11'd517 : tab = 23'b10011000101110001101000;
11'd518 : tab = 23'b10011000100100000000110;
11'd519 : tab = 23'b10011000011001110101000;
11'd520 : tab = 23'b10011000001111101001100;
11'd521 : tab = 23'b10011000000101011110110;
11'd522 : tab = 23'b10010111111011010100100;
11'd523 : tab = 23'b10010111110001001010110;
11'd524 : tab = 23'b10010111100111000001100;
11'd525 : tab = 23'b10010111011100111000110;
11'd526 : tab = 23'b10010111010010110000100;
11'd527 : tab = 23'b10010111001000101000110;
11'd528 : tab = 23'b10010110111110100001100;
11'd529 : tab = 23'b10010110110100011010110;
11'd530 : tab = 23'b10010110101010010100100;
11'd531 : tab = 23'b10010110100000001110110;
11'd532 : tab = 23'b10010110010110001001100;
11'd533 : tab = 23'b10010110001100000100110;
11'd534 : tab = 23'b10010110000010000000101;
11'd535 : tab = 23'b10010101110111111100111;
11'd536 : tab = 23'b10010101101101111001101;
11'd537 : tab = 23'b10010101100011110110111;
11'd538 : tab = 23'b10010101011001110100101;
11'd539 : tab = 23'b10010101001111110010111;
11'd540 : tab = 23'b10010101000101110001101;
11'd541 : tab = 23'b10010100111011110000111;
11'd542 : tab = 23'b10010100110001110000100;
11'd543 : tab = 23'b10010100100111110000110;
11'd544 : tab = 23'b10010100011101110001100;
11'd545 : tab = 23'b10010100010011110010110;
11'd546 : tab = 23'b10010100001001110100100;
11'd547 : tab = 23'b10010011111111110110110;
11'd548 : tab = 23'b10010011110101111001011;
11'd549 : tab = 23'b10010011101011111100100;
11'd550 : tab = 23'b10010011100010000000010;
11'd551 : tab = 23'b10010011011000000100011;
11'd552 : tab = 23'b10010011001110001001000;
11'd553 : tab = 23'b10010011000100001110001;
11'd554 : tab = 23'b10010010111010010011110;
11'd555 : tab = 23'b10010010110000011001111;
11'd556 : tab = 23'b10010010100110100000100;
11'd557 : tab = 23'b10010010011100100111101;
11'd558 : tab = 23'b10010010010010101111001;
11'd559 : tab = 23'b10010010001000110111010;
11'd560 : tab = 23'b10010001111110111111110;
11'd561 : tab = 23'b10010001110101001000110;
11'd562 : tab = 23'b10010001101011010010010;
11'd563 : tab = 23'b10010001100001011100010;
11'd564 : tab = 23'b10010001010111100110110;
11'd565 : tab = 23'b10010001001101110001110;
11'd566 : tab = 23'b10010001000011111101010;
11'd567 : tab = 23'b10010000111010001001000;
11'd568 : tab = 23'b10010000110000010101100;
11'd569 : tab = 23'b10010000100110100010011;
11'd570 : tab = 23'b10010000011100101111110;
11'd571 : tab = 23'b10010000010010111101100;
11'd572 : tab = 23'b10010000001001001011111;
11'd573 : tab = 23'b10001111111111011010101;
11'd574 : tab = 23'b10001111110101101010000;
11'd575 : tab = 23'b10001111101011111001110;
11'd576 : tab = 23'b10001111100010001001110;
11'd577 : tab = 23'b10001111011000011010100;
11'd578 : tab = 23'b10001111001110101011110;
11'd579 : tab = 23'b10001111000100111101011;
11'd580 : tab = 23'b10001110111011001111100;
11'd581 : tab = 23'b10001110110001100010001;
11'd582 : tab = 23'b10001110100111110101001;
11'd583 : tab = 23'b10001110011110001000110;
11'd584 : tab = 23'b10001110010100011100110;
11'd585 : tab = 23'b10001110001010110001010;
11'd586 : tab = 23'b10001110000001000110000;
11'd587 : tab = 23'b10001101110111011011100;
11'd588 : tab = 23'b10001101101101110001011;
11'd589 : tab = 23'b10001101100100000111110;
11'd590 : tab = 23'b10001101011010011110100;
11'd591 : tab = 23'b10001101010000110101111;
11'd592 : tab = 23'b10001101000111001101101;
11'd593 : tab = 23'b10001100111101100101110;
11'd594 : tab = 23'b10001100110011111110100;
11'd595 : tab = 23'b10001100101010010111110;
11'd596 : tab = 23'b10001100100000110001010;
11'd597 : tab = 23'b10001100010111001011011;
11'd598 : tab = 23'b10001100001101100110000;
11'd599 : tab = 23'b10001100000100000001000;
11'd600 : tab = 23'b10001011111010011100100;
11'd601 : tab = 23'b10001011110000111000011;
11'd602 : tab = 23'b10001011100111010100110;
11'd603 : tab = 23'b10001011011101110001101;
11'd604 : tab = 23'b10001011010100001111000;
11'd605 : tab = 23'b10001011001010101100110;
11'd606 : tab = 23'b10001011000001001011000;
11'd607 : tab = 23'b10001010110111101001110;
11'd608 : tab = 23'b10001010101110001000110;
11'd609 : tab = 23'b10001010100100101000100;
11'd610 : tab = 23'b10001010011011001000100;
11'd611 : tab = 23'b10001010010001101001000;
11'd612 : tab = 23'b10001010001000001010000;
11'd613 : tab = 23'b10001001111110101011100;
11'd614 : tab = 23'b10001001110101001101011;
11'd615 : tab = 23'b10001001101011101111110;
11'd616 : tab = 23'b10001001100010010010100;
11'd617 : tab = 23'b10001001011000110101110;
11'd618 : tab = 23'b10001001001111011001100;
11'd619 : tab = 23'b10001001000101111101110;
11'd620 : tab = 23'b10001000111100100010011;
11'd621 : tab = 23'b10001000110011000111011;
11'd622 : tab = 23'b10001000101001101101000;
11'd623 : tab = 23'b10001000100000010011000;
11'd624 : tab = 23'b10001000010110111001011;
11'd625 : tab = 23'b10001000001101100000010;
11'd626 : tab = 23'b10001000000100000111100;
11'd627 : tab = 23'b10000111111010101111010;
11'd628 : tab = 23'b10000111110001010111100;
11'd629 : tab = 23'b10000111101000000000010;
11'd630 : tab = 23'b10000111011110101001011;
11'd631 : tab = 23'b10000111010101010011000;
11'd632 : tab = 23'b10000111001011111101000;
11'd633 : tab = 23'b10000111000010100111011;
11'd634 : tab = 23'b10000110111001010010010;
11'd635 : tab = 23'b10000110101111111101101;
11'd636 : tab = 23'b10000110100110101001100;
11'd637 : tab = 23'b10000110011101010101110;
11'd638 : tab = 23'b10000110010100000010011;
11'd639 : tab = 23'b10000110001010101111100;
11'd640 : tab = 23'b10000110000001011101000;
11'd641 : tab = 23'b10000101111000001011000;
11'd642 : tab = 23'b10000101101110111001100;
11'd643 : tab = 23'b10000101100101101000011;
11'd644 : tab = 23'b10000101011100010111110;
11'd645 : tab = 23'b10000101010011000111100;
11'd646 : tab = 23'b10000101001001110111110;
11'd647 : tab = 23'b10000101000000101000011;
11'd648 : tab = 23'b10000100110111011001100;
11'd649 : tab = 23'b10000100101110001011000;
11'd650 : tab = 23'b10000100100100111101000;
11'd651 : tab = 23'b10000100011011101111011;
11'd652 : tab = 23'b10000100010010100010010;
11'd653 : tab = 23'b10000100001001010101100;
11'd654 : tab = 23'b10000100000000001001010;
11'd655 : tab = 23'b10000011110110111101011;
11'd656 : tab = 23'b10000011101101110010000;
11'd657 : tab = 23'b10000011100100100111000;
11'd658 : tab = 23'b10000011011011011100100;
11'd659 : tab = 23'b10000011010010010010010;
11'd660 : tab = 23'b10000011001001001000101;
11'd661 : tab = 23'b10000010111111111111011;
11'd662 : tab = 23'b10000010110110110110100;
11'd663 : tab = 23'b10000010101101101110001;
11'd664 : tab = 23'b10000010100100100110010;
11'd665 : tab = 23'b10000010011011011110110;
11'd666 : tab = 23'b10000010010010010111101;
11'd667 : tab = 23'b10000010001001010001000;
11'd668 : tab = 23'b10000010000000001010110;
11'd669 : tab = 23'b10000001110111000100111;
11'd670 : tab = 23'b10000001101101111111100;
11'd671 : tab = 23'b10000001100100111010100;
11'd672 : tab = 23'b10000001011011110110000;
11'd673 : tab = 23'b10000001010010110001111;
11'd674 : tab = 23'b10000001001001101110010;
11'd675 : tab = 23'b10000001000000101011000;
11'd676 : tab = 23'b10000000110111101000001;
11'd677 : tab = 23'b10000000101110100101110;
11'd678 : tab = 23'b10000000100101100011110;
11'd679 : tab = 23'b10000000011100100010010;
11'd680 : tab = 23'b10000000010011100001001;
11'd681 : tab = 23'b10000000001010100000100;
11'd682 : tab = 23'b10000000000001100000001;
11'd683 : tab = 23'b01111111111000100000010;
11'd684 : tab = 23'b01111111101111100000110;
11'd685 : tab = 23'b01111111100110100001110;
11'd686 : tab = 23'b01111111011101100011010;
11'd687 : tab = 23'b01111111010100100101000;
11'd688 : tab = 23'b01111111001011100111010;
11'd689 : tab = 23'b01111111000010101010000;
11'd690 : tab = 23'b01111110111001101101000;
11'd691 : tab = 23'b01111110110000110000100;
11'd692 : tab = 23'b01111110100111110100100;
11'd693 : tab = 23'b01111110011110111000110;
11'd694 : tab = 23'b01111110010101111101100;
11'd695 : tab = 23'b01111110001101000010110;
11'd696 : tab = 23'b01111110000100001000010;
11'd697 : tab = 23'b01111101111011001110010;
11'd698 : tab = 23'b01111101110010010100110;
11'd699 : tab = 23'b01111101101001011011100;
11'd700 : tab = 23'b01111101100000100010110;
11'd701 : tab = 23'b01111101010111101010011;
11'd702 : tab = 23'b01111101001110110010100;
11'd703 : tab = 23'b01111101000101111011000;
11'd704 : tab = 23'b01111100111101000011111;
11'd705 : tab = 23'b01111100110100001101010;
11'd706 : tab = 23'b01111100101011010110111;
11'd707 : tab = 23'b01111100100010100001000;
11'd708 : tab = 23'b01111100011001101011100;
11'd709 : tab = 23'b01111100010000110110100;
11'd710 : tab = 23'b01111100001000000001111;
11'd711 : tab = 23'b01111011111111001101110;
11'd712 : tab = 23'b01111011110110011001111;
11'd713 : tab = 23'b01111011101101100110100;
11'd714 : tab = 23'b01111011100100110011100;
11'd715 : tab = 23'b01111011011100000000110;
11'd716 : tab = 23'b01111011010011001110101;
11'd717 : tab = 23'b01111011001010011100110;
11'd718 : tab = 23'b01111011000001101011100;
11'd719 : tab = 23'b01111010111000111010100;
11'd720 : tab = 23'b01111010110000001001111;
11'd721 : tab = 23'b01111010100111011001110;
11'd722 : tab = 23'b01111010011110101010000;
11'd723 : tab = 23'b01111010010101111010101;
11'd724 : tab = 23'b01111010001101001011110;
11'd725 : tab = 23'b01111010000100011101001;
11'd726 : tab = 23'b01111001111011101111000;
11'd727 : tab = 23'b01111001110011000001010;
11'd728 : tab = 23'b01111001101010010011111;
11'd729 : tab = 23'b01111001100001100111000;
11'd730 : tab = 23'b01111001011000111010100;
11'd731 : tab = 23'b01111001010000001110010;
11'd732 : tab = 23'b01111001000111100010100;
11'd733 : tab = 23'b01111000111110110111010;
11'd734 : tab = 23'b01111000110110001100010;
11'd735 : tab = 23'b01111000101101100001110;
11'd736 : tab = 23'b01111000100100110111101;
11'd737 : tab = 23'b01111000011100001101110;
11'd738 : tab = 23'b01111000010011100100100;
11'd739 : tab = 23'b01111000001010111011100;
11'd740 : tab = 23'b01111000000010010011000;
11'd741 : tab = 23'b01110111111001101010110;
11'd742 : tab = 23'b01110111110001000011000;
11'd743 : tab = 23'b01110111101000011011110;
11'd744 : tab = 23'b01110111011111110100110;
11'd745 : tab = 23'b01110111010111001110001;
11'd746 : tab = 23'b01110111001110101000000;
11'd747 : tab = 23'b01110111000110000010010;
11'd748 : tab = 23'b01110110111101011100110;
11'd749 : tab = 23'b01110110110100110111110;
11'd750 : tab = 23'b01110110101100010011010;
11'd751 : tab = 23'b01110110100011101111000;
11'd752 : tab = 23'b01110110011011001011001;
11'd753 : tab = 23'b01110110010010100111110;
11'd754 : tab = 23'b01110110001010000100101;
11'd755 : tab = 23'b01110110000001100010000;
11'd756 : tab = 23'b01110101111000111111110;
11'd757 : tab = 23'b01110101110000011101111;
11'd758 : tab = 23'b01110101100111111100011;
11'd759 : tab = 23'b01110101011111011011010;
11'd760 : tab = 23'b01110101010110111010100;
11'd761 : tab = 23'b01110101001110011010010;
11'd762 : tab = 23'b01110101000101111010010;
11'd763 : tab = 23'b01110100111101011010110;
11'd764 : tab = 23'b01110100110100111011100;
11'd765 : tab = 23'b01110100101100011100110;
11'd766 : tab = 23'b01110100100011111110100;
11'd767 : tab = 23'b01110100011011100000100;
11'd768 : tab = 23'b01110100010011000010110;
11'd769 : tab = 23'b01110100001010100101100;
11'd770 : tab = 23'b01110100000010001000110;
11'd771 : tab = 23'b01110011111001101100010;
11'd772 : tab = 23'b01110011110001010000001;
11'd773 : tab = 23'b01110011101000110100100;
11'd774 : tab = 23'b01110011100000011001001;
11'd775 : tab = 23'b01110011010111111110010;
11'd776 : tab = 23'b01110011001111100011101;
11'd777 : tab = 23'b01110011000111001001100;
11'd778 : tab = 23'b01110010111110101111110;
11'd779 : tab = 23'b01110010110110010110010;
11'd780 : tab = 23'b01110010101101111101010;
11'd781 : tab = 23'b01110010100101100100100;
11'd782 : tab = 23'b01110010011101001100010;
11'd783 : tab = 23'b01110010010100110100100;
11'd784 : tab = 23'b01110010001100011100111;
11'd785 : tab = 23'b01110010000100000101110;
11'd786 : tab = 23'b01110001111011101111000;
11'd787 : tab = 23'b01110001110011011000101;
11'd788 : tab = 23'b01110001101011000010101;
11'd789 : tab = 23'b01110001100010101101000;
11'd790 : tab = 23'b01110001011010010111110;
11'd791 : tab = 23'b01110001010010000010110;
11'd792 : tab = 23'b01110001001001101110010;
11'd793 : tab = 23'b01110001000001011010010;
11'd794 : tab = 23'b01110000111001000110100;
11'd795 : tab = 23'b01110000110000110011000;
11'd796 : tab = 23'b01110000101000100000000;
11'd797 : tab = 23'b01110000100000001101100;
11'd798 : tab = 23'b01110000010111111011010;
11'd799 : tab = 23'b01110000001111101001010;
11'd800 : tab = 23'b01110000000111010111110;
11'd801 : tab = 23'b01101111111111000110101;
11'd802 : tab = 23'b01101111110110110101111;
11'd803 : tab = 23'b01101111101110100101100;
11'd804 : tab = 23'b01101111100110010101011;
11'd805 : tab = 23'b01101111011110000101110;
11'd806 : tab = 23'b01101111010101110110100;
11'd807 : tab = 23'b01101111001101100111100;
11'd808 : tab = 23'b01101111000101011001000;
11'd809 : tab = 23'b01101110111101001010110;
11'd810 : tab = 23'b01101110110100111101000;
11'd811 : tab = 23'b01101110101100101111100;
11'd812 : tab = 23'b01101110100100100010100;
11'd813 : tab = 23'b01101110011100010101110;
11'd814 : tab = 23'b01101110010100001001011;
11'd815 : tab = 23'b01101110001011111101011;
11'd816 : tab = 23'b01101110000011110001110;
11'd817 : tab = 23'b01101101111011100110100;
11'd818 : tab = 23'b01101101110011011011101;
11'd819 : tab = 23'b01101101101011010001001;
11'd820 : tab = 23'b01101101100011000111000;
11'd821 : tab = 23'b01101101011010111101001;
11'd822 : tab = 23'b01101101010010110011110;
11'd823 : tab = 23'b01101101001010101010101;
11'd824 : tab = 23'b01101101000010100010000;
11'd825 : tab = 23'b01101100111010011001101;
11'd826 : tab = 23'b01101100110010010001101;
11'd827 : tab = 23'b01101100101010001010000;
11'd828 : tab = 23'b01101100100010000010110;
11'd829 : tab = 23'b01101100011001111011111;
11'd830 : tab = 23'b01101100010001110101011;
11'd831 : tab = 23'b01101100001001101111010;
11'd832 : tab = 23'b01101100000001101001011;
11'd833 : tab = 23'b01101011111001100011111;
11'd834 : tab = 23'b01101011110001011110110;
11'd835 : tab = 23'b01101011101001011010000;
11'd836 : tab = 23'b01101011100001010101110;
11'd837 : tab = 23'b01101011011001010001101;
11'd838 : tab = 23'b01101011010001001110000;
11'd839 : tab = 23'b01101011001001001010101;
11'd840 : tab = 23'b01101011000001000111110;
11'd841 : tab = 23'b01101010111001000101001;
11'd842 : tab = 23'b01101010110001000010111;
11'd843 : tab = 23'b01101010101001000001000;
11'd844 : tab = 23'b01101010100000111111100;
11'd845 : tab = 23'b01101010011000111110010;
11'd846 : tab = 23'b01101010010000111101100;
11'd847 : tab = 23'b01101010001000111101000;
11'd848 : tab = 23'b01101010000000111101000;
11'd849 : tab = 23'b01101001111000111101001;
11'd850 : tab = 23'b01101001110000111101110;
11'd851 : tab = 23'b01101001101000111110110;
11'd852 : tab = 23'b01101001100001000000000;
11'd853 : tab = 23'b01101001011001000001101;
11'd854 : tab = 23'b01101001010001000011110;
11'd855 : tab = 23'b01101001001001000110000;
11'd856 : tab = 23'b01101001000001001000110;
11'd857 : tab = 23'b01101000111001001011110;
11'd858 : tab = 23'b01101000110001001111010;
11'd859 : tab = 23'b01101000101001010011000;
11'd860 : tab = 23'b01101000100001010111000;
11'd861 : tab = 23'b01101000011001011011100;
11'd862 : tab = 23'b01101000010001100000010;
11'd863 : tab = 23'b01101000001001100101100;
11'd864 : tab = 23'b01101000000001101011000;
11'd865 : tab = 23'b01100111111001110000110;
11'd866 : tab = 23'b01100111110001110111000;
11'd867 : tab = 23'b01100111101001111101100;
11'd868 : tab = 23'b01100111100010000100100;
11'd869 : tab = 23'b01100111011010001011110;
11'd870 : tab = 23'b01100111010010010011010;
11'd871 : tab = 23'b01100111001010011011010;
11'd872 : tab = 23'b01100111000010100011100;
11'd873 : tab = 23'b01100110111010101100001;
11'd874 : tab = 23'b01100110110010110101001;
11'd875 : tab = 23'b01100110101010111110011;
11'd876 : tab = 23'b01100110100011001000000;
11'd877 : tab = 23'b01100110011011010010000;
11'd878 : tab = 23'b01100110010011011100010;
11'd879 : tab = 23'b01100110001011100111000;
11'd880 : tab = 23'b01100110000011110010000;
11'd881 : tab = 23'b01100101111011111101100;
11'd882 : tab = 23'b01100101110100001001001;
11'd883 : tab = 23'b01100101101100010101010;
11'd884 : tab = 23'b01100101100100100001100;
11'd885 : tab = 23'b01100101011100101110010;
11'd886 : tab = 23'b01100101010100111011011;
11'd887 : tab = 23'b01100101001101001000110;
11'd888 : tab = 23'b01100101000101010110100;
11'd889 : tab = 23'b01100100111101100100110;
11'd890 : tab = 23'b01100100110101110011000;
11'd891 : tab = 23'b01100100101110000001110;
11'd892 : tab = 23'b01100100100110010001000;
11'd893 : tab = 23'b01100100011110100000011;
11'd894 : tab = 23'b01100100010110110000001;
11'd895 : tab = 23'b01100100001111000000010;
11'd896 : tab = 23'b01100100000111010000110;
11'd897 : tab = 23'b01100011111111100001100;
11'd898 : tab = 23'b01100011110111110010101;
11'd899 : tab = 23'b01100011110000000100001;
11'd900 : tab = 23'b01100011101000010110000;
11'd901 : tab = 23'b01100011100000101000000;
11'd902 : tab = 23'b01100011011000111010100;
11'd903 : tab = 23'b01100011010001001101010;
11'd904 : tab = 23'b01100011001001100000100;
11'd905 : tab = 23'b01100011000001110011111;
11'd906 : tab = 23'b01100010111010000111110;
11'd907 : tab = 23'b01100010110010011011110;
11'd908 : tab = 23'b01100010101010110000010;
11'd909 : tab = 23'b01100010100011000101001;
11'd910 : tab = 23'b01100010011011011010010;
11'd911 : tab = 23'b01100010010011101111110;
11'd912 : tab = 23'b01100010001100000101100;
11'd913 : tab = 23'b01100010000100011011101;
11'd914 : tab = 23'b01100001111100110010001;
11'd915 : tab = 23'b01100001110101001000111;
11'd916 : tab = 23'b01100001101101100000000;
11'd917 : tab = 23'b01100001100101110111100;
11'd918 : tab = 23'b01100001011110001111010;
11'd919 : tab = 23'b01100001010110100111010;
11'd920 : tab = 23'b01100001001110111111110;
11'd921 : tab = 23'b01100001000111011000100;
11'd922 : tab = 23'b01100000111111110001100;
11'd923 : tab = 23'b01100000111000001011000;
11'd924 : tab = 23'b01100000110000100100110;
11'd925 : tab = 23'b01100000101000111110110;
11'd926 : tab = 23'b01100000100001011001010;
11'd927 : tab = 23'b01100000011001110100000;
11'd928 : tab = 23'b01100000010010001111000;
11'd929 : tab = 23'b01100000001010101010100;
11'd930 : tab = 23'b01100000000011000110001;
11'd931 : tab = 23'b01011111111011100010001;
11'd932 : tab = 23'b01011111110011111110100;
11'd933 : tab = 23'b01011111101100011011010;
11'd934 : tab = 23'b01011111100100111000010;
11'd935 : tab = 23'b01011111011101010101100;
11'd936 : tab = 23'b01011111010101110011010;
11'd937 : tab = 23'b01011111001110010001001;
11'd938 : tab = 23'b01011111000110101111100;
11'd939 : tab = 23'b01011110111111001110000;
11'd940 : tab = 23'b01011110110111101101000;
11'd941 : tab = 23'b01011110110000001100010;
11'd942 : tab = 23'b01011110101000101011110;
11'd943 : tab = 23'b01011110100001001011110;
11'd944 : tab = 23'b01011110011001101100000;
11'd945 : tab = 23'b01011110010010001100100;
11'd946 : tab = 23'b01011110001010101101100;
11'd947 : tab = 23'b01011110000011001110100;
11'd948 : tab = 23'b01011101111011110000001;
11'd949 : tab = 23'b01011101110100010010000;
11'd950 : tab = 23'b01011101101100110100000;
11'd951 : tab = 23'b01011101100101010110100;
11'd952 : tab = 23'b01011101011101111001010;
11'd953 : tab = 23'b01011101010110011100100;
11'd954 : tab = 23'b01011101001110111111110;
11'd955 : tab = 23'b01011101000111100011100;
11'd956 : tab = 23'b01011101000000000111100;
11'd957 : tab = 23'b01011100111000101100000;
11'd958 : tab = 23'b01011100110001010000101;
11'd959 : tab = 23'b01011100101001110101101;
11'd960 : tab = 23'b01011100100010011011000;
11'd961 : tab = 23'b01011100011011000000100;
11'd962 : tab = 23'b01011100010011100110100;
11'd963 : tab = 23'b01011100001100001100110;
11'd964 : tab = 23'b01011100000100110011011;
11'd965 : tab = 23'b01011011111101011010010;
11'd966 : tab = 23'b01011011110110000001100;
11'd967 : tab = 23'b01011011101110101001000;
11'd968 : tab = 23'b01011011100111010000110;
11'd969 : tab = 23'b01011011011111111001000;
11'd970 : tab = 23'b01011011011000100001100;
11'd971 : tab = 23'b01011011010001001010010;
11'd972 : tab = 23'b01011011001001110011010;
11'd973 : tab = 23'b01011011000010011100110;
11'd974 : tab = 23'b01011010111011000110011;
11'd975 : tab = 23'b01011010110011110000011;
11'd976 : tab = 23'b01011010101100011010110;
11'd977 : tab = 23'b01011010100101000101010;
11'd978 : tab = 23'b01011010011101110000010;
11'd979 : tab = 23'b01011010010110011011100;
11'd980 : tab = 23'b01011010001111000111001;
11'd981 : tab = 23'b01011010000111110011000;
11'd982 : tab = 23'b01011010000000011111010;
11'd983 : tab = 23'b01011001111001001011101;
11'd984 : tab = 23'b01011001110001111000100;
11'd985 : tab = 23'b01011001101010100101100;
11'd986 : tab = 23'b01011001100011010011000;
11'd987 : tab = 23'b01011001011100000000110;
11'd988 : tab = 23'b01011001010100101110110;
11'd989 : tab = 23'b01011001001101011101000;
11'd990 : tab = 23'b01011001000110001011110;
11'd991 : tab = 23'b01011000111110111010110;
11'd992 : tab = 23'b01011000110111101010000;
11'd993 : tab = 23'b01011000110000011001100;
11'd994 : tab = 23'b01011000101001001001100;
11'd995 : tab = 23'b01011000100001111001100;
11'd996 : tab = 23'b01011000011010101010000;
11'd997 : tab = 23'b01011000010011011010110;
11'd998 : tab = 23'b01011000001100001100000;
11'd999 : tab = 23'b01011000000100111101010;
11'd1000 : tab = 23'b01010111111101101111000;
11'd1001 : tab = 23'b01010111110110100001000;
11'd1002 : tab = 23'b01010111101111010011010;
11'd1003 : tab = 23'b01010111101000000110000;
11'd1004 : tab = 23'b01010111100000111000110;
11'd1005 : tab = 23'b01010111011001101100000;
11'd1006 : tab = 23'b01010111010010011111100;
11'd1007 : tab = 23'b01010111001011010011010;
11'd1008 : tab = 23'b01010111000100000111100;
11'd1009 : tab = 23'b01010110111100111011110;
11'd1010 : tab = 23'b01010110110101110000100;
11'd1011 : tab = 23'b01010110101110100101100;
11'd1012 : tab = 23'b01010110100111011010111;
11'd1013 : tab = 23'b01010110100000010000100;
11'd1014 : tab = 23'b01010110011001000110011;
11'd1015 : tab = 23'b01010110010001111100101;
11'd1016 : tab = 23'b01010110001010110011001;
11'd1017 : tab = 23'b01010110000011101010000;
11'd1018 : tab = 23'b01010101111100100001000;
11'd1019 : tab = 23'b01010101110101011000100;
11'd1020 : tab = 23'b01010101101110010000001;
11'd1021 : tab = 23'b01010101100111001000001;
11'd1022 : tab = 23'b01010101100000000000100;
11'd1023 : tab = 23'b01010101011000111001000;
11'd1024 : tab = 23'b01010101010001110010000;
11'd1025 : tab = 23'b01010101001010101011001;
11'd1026 : tab = 23'b01010101000011100100101;
11'd1027 : tab = 23'b01010100111100011110011;
11'd1028 : tab = 23'b01010100110101011000100;
11'd1029 : tab = 23'b01010100101110010010110;
11'd1030 : tab = 23'b01010100100111001101100;
11'd1031 : tab = 23'b01010100100000001000011;
11'd1032 : tab = 23'b01010100011001000011101;
11'd1033 : tab = 23'b01010100010001111111010;
11'd1034 : tab = 23'b01010100001010111011000;
11'd1035 : tab = 23'b01010100000011110111010;
11'd1036 : tab = 23'b01010011111100110011100;
11'd1037 : tab = 23'b01010011110101110000010;
11'd1038 : tab = 23'b01010011101110101101010;
11'd1039 : tab = 23'b01010011100111101010101;
11'd1040 : tab = 23'b01010011100000101000010;
11'd1041 : tab = 23'b01010011011001100110000;
11'd1042 : tab = 23'b01010011010010100100010;
11'd1043 : tab = 23'b01010011001011100010110;
11'd1044 : tab = 23'b01010011000100100001100;
11'd1045 : tab = 23'b01010010111101100000100;
11'd1046 : tab = 23'b01010010110110011111111;
11'd1047 : tab = 23'b01010010101111011111100;
11'd1048 : tab = 23'b01010010101000011111100;
11'd1049 : tab = 23'b01010010100001011111101;
11'd1050 : tab = 23'b01010010011010100000001;
11'd1051 : tab = 23'b01010010010011100000111;
11'd1052 : tab = 23'b01010010001100100010000;
11'd1053 : tab = 23'b01010010000101100011010;
11'd1054 : tab = 23'b01010001111110100101000;
11'd1055 : tab = 23'b01010001110111100111000;
11'd1056 : tab = 23'b01010001110000101001001;
11'd1057 : tab = 23'b01010001101001101011101;
11'd1058 : tab = 23'b01010001100010101110100;
11'd1059 : tab = 23'b01010001011011110001100;
11'd1060 : tab = 23'b01010001010100110101000;
11'd1061 : tab = 23'b01010001001101111000100;
11'd1062 : tab = 23'b01010001000110111100100;
11'd1063 : tab = 23'b01010001000000000000110;
11'd1064 : tab = 23'b01010000111001000101010;
11'd1065 : tab = 23'b01010000110010001010000;
11'd1066 : tab = 23'b01010000101011001111001;
11'd1067 : tab = 23'b01010000100100010100100;
11'd1068 : tab = 23'b01010000011101011010010;
11'd1069 : tab = 23'b01010000010110100000000;
11'd1070 : tab = 23'b01010000001111100110010;
11'd1071 : tab = 23'b01010000001000101100111;
11'd1072 : tab = 23'b01010000000001110011101;
11'd1073 : tab = 23'b01001111111010111010110;
11'd1074 : tab = 23'b01001111110100000010000;
11'd1075 : tab = 23'b01001111101101001001110;
11'd1076 : tab = 23'b01001111100110010001100;
11'd1077 : tab = 23'b01001111011111011001110;
11'd1078 : tab = 23'b01001111011000100010010;
11'd1079 : tab = 23'b01001111010001101011000;
11'd1080 : tab = 23'b01001111001010110100000;
11'd1081 : tab = 23'b01001111000011111101011;
11'd1082 : tab = 23'b01001110111101000111000;
11'd1083 : tab = 23'b01001110110110010000110;
11'd1084 : tab = 23'b01001110101111011011000;
11'd1085 : tab = 23'b01001110101000100101100;
11'd1086 : tab = 23'b01001110100001110000001;
11'd1087 : tab = 23'b01001110011010111011001;
11'd1088 : tab = 23'b01001110010100000110011;
11'd1089 : tab = 23'b01001110001101010010000;
11'd1090 : tab = 23'b01001110000110011101110;
11'd1091 : tab = 23'b01001101111111101010000;
11'd1092 : tab = 23'b01001101111000110110010;
11'd1093 : tab = 23'b01001101110010000011000;
11'd1094 : tab = 23'b01001101101011001111111;
11'd1095 : tab = 23'b01001101100100011101001;
11'd1096 : tab = 23'b01001101011101101010101;
11'd1097 : tab = 23'b01001101010110111000011;
11'd1098 : tab = 23'b01001101010000000110100;
11'd1099 : tab = 23'b01001101001001010100110;
11'd1100 : tab = 23'b01001101000010100011010;
11'd1101 : tab = 23'b01001100111011110010010;
11'd1102 : tab = 23'b01001100110101000001011;
11'd1103 : tab = 23'b01001100101110010000110;
11'd1104 : tab = 23'b01001100100111100000100;
11'd1105 : tab = 23'b01001100100000110000100;
11'd1106 : tab = 23'b01001100011010000000110;
11'd1107 : tab = 23'b01001100010011010001010;
11'd1108 : tab = 23'b01001100001100100010000;
11'd1109 : tab = 23'b01001100000101110011001;
11'd1110 : tab = 23'b01001011111111000100100;
11'd1111 : tab = 23'b01001011111000010110000;
11'd1112 : tab = 23'b01001011110001101000000;
11'd1113 : tab = 23'b01001011101010111010000;
11'd1114 : tab = 23'b01001011100100001100100;
11'd1115 : tab = 23'b01001011011101011111010;
11'd1116 : tab = 23'b01001011010110110010010;
11'd1117 : tab = 23'b01001011010000000101011;
11'd1118 : tab = 23'b01001011001001011000111;
11'd1119 : tab = 23'b01001011000010101100110;
11'd1120 : tab = 23'b01001010111100000000110;
11'd1121 : tab = 23'b01001010110101010101001;
11'd1122 : tab = 23'b01001010101110101001110;
11'd1123 : tab = 23'b01001010100111111110100;
11'd1124 : tab = 23'b01001010100001010011110;
11'd1125 : tab = 23'b01001010011010101001000;
11'd1126 : tab = 23'b01001010010011111110110;
11'd1127 : tab = 23'b01001010001101010100110;
11'd1128 : tab = 23'b01001010000110101010111;
11'd1129 : tab = 23'b01001010000000000001011;
11'd1130 : tab = 23'b01001001111001011000001;
11'd1131 : tab = 23'b01001001110010101111001;
11'd1132 : tab = 23'b01001001101100000110011;
11'd1133 : tab = 23'b01001001100101011110000;
11'd1134 : tab = 23'b01001001011110110101110;
11'd1135 : tab = 23'b01001001011000001101110;
11'd1136 : tab = 23'b01001001010001100110010;
11'd1137 : tab = 23'b01001001001010111110110;
11'd1138 : tab = 23'b01001001000100010111110;
11'd1139 : tab = 23'b01001000111101110000110;
11'd1140 : tab = 23'b01001000110111001010010;
11'd1141 : tab = 23'b01001000110000100011111;
11'd1142 : tab = 23'b01001000101001111101110;
11'd1143 : tab = 23'b01001000100011011000000;
11'd1144 : tab = 23'b01001000011100110010100;
11'd1145 : tab = 23'b01001000010110001101010;
11'd1146 : tab = 23'b01001000001111101000010;
11'd1147 : tab = 23'b01001000001001000011100;
11'd1148 : tab = 23'b01001000000010011111000;
11'd1149 : tab = 23'b01000111111011111010110;
11'd1150 : tab = 23'b01000111110101010110110;
11'd1151 : tab = 23'b01000111101110110011001;
11'd1152 : tab = 23'b01000111101000001111110;
11'd1153 : tab = 23'b01000111100001101100100;
11'd1154 : tab = 23'b01000111011011001001101;
11'd1155 : tab = 23'b01000111010100100111000;
11'd1156 : tab = 23'b01000111001110000100100;
11'd1157 : tab = 23'b01000111000111100010100;
11'd1158 : tab = 23'b01000111000001000000100;
11'd1159 : tab = 23'b01000110111010011111000;
11'd1160 : tab = 23'b01000110110011111101110;
11'd1161 : tab = 23'b01000110101101011100100;
11'd1162 : tab = 23'b01000110100110111011110;
11'd1163 : tab = 23'b01000110100000011011010;
11'd1164 : tab = 23'b01000110011001111010111;
11'd1165 : tab = 23'b01000110010011011010110;
11'd1166 : tab = 23'b01000110001100111011000;
11'd1167 : tab = 23'b01000110000110011011100;
11'd1168 : tab = 23'b01000101111111111100010;
11'd1169 : tab = 23'b01000101111001011101010;
11'd1170 : tab = 23'b01000101110010111110100;
11'd1171 : tab = 23'b01000101101100100000000;
11'd1172 : tab = 23'b01000101100110000001110;
11'd1173 : tab = 23'b01000101011111100011110;
11'd1174 : tab = 23'b01000101011001000110001;
11'd1175 : tab = 23'b01000101010010101000101;
11'd1176 : tab = 23'b01000101001100001011011;
11'd1177 : tab = 23'b01000101000101101110100;
11'd1178 : tab = 23'b01000100111111010001110;
11'd1179 : tab = 23'b01000100111000110101010;
11'd1180 : tab = 23'b01000100110010011001001;
11'd1181 : tab = 23'b01000100101011111101010;
11'd1182 : tab = 23'b01000100100101100001100;
11'd1183 : tab = 23'b01000100011111000110001;
11'd1184 : tab = 23'b01000100011000101011000;
11'd1185 : tab = 23'b01000100010010010000000;
11'd1186 : tab = 23'b01000100001011110101011;
11'd1187 : tab = 23'b01000100000101011011000;
11'd1188 : tab = 23'b01000011111111000000110;
11'd1189 : tab = 23'b01000011111000100111000;
11'd1190 : tab = 23'b01000011110010001101010;
11'd1191 : tab = 23'b01000011101011110011111;
11'd1192 : tab = 23'b01000011100101011010110;
11'd1193 : tab = 23'b01000011011111000001110;
11'd1194 : tab = 23'b01000011011000101001010;
11'd1195 : tab = 23'b01000011010010010000110;
11'd1196 : tab = 23'b01000011001011111000110;
11'd1197 : tab = 23'b01000011000101100000110;
11'd1198 : tab = 23'b01000010111111001001010;
11'd1199 : tab = 23'b01000010111000110001110;
11'd1200 : tab = 23'b01000010110010011010110;
11'd1201 : tab = 23'b01000010101100000011110;
11'd1202 : tab = 23'b01000010100101101101010;
11'd1203 : tab = 23'b01000010011111010110110;
11'd1204 : tab = 23'b01000010011001000000110;
11'd1205 : tab = 23'b01000010010010101010110;
11'd1206 : tab = 23'b01000010001100010101010;
11'd1207 : tab = 23'b01000010000101111111110;
11'd1208 : tab = 23'b01000001111111101010110;
11'd1209 : tab = 23'b01000001111001010101110;
11'd1210 : tab = 23'b01000001110011000001010;
11'd1211 : tab = 23'b01000001101100101100110;
11'd1212 : tab = 23'b01000001100110011000110;
11'd1213 : tab = 23'b01000001100000000100110;
11'd1214 : tab = 23'b01000001011001110001010;
11'd1215 : tab = 23'b01000001010011011101110;
11'd1216 : tab = 23'b01000001001101001010101;
11'd1217 : tab = 23'b01000001000110110111110;
11'd1218 : tab = 23'b01000001000000100101000;
11'd1219 : tab = 23'b01000000111010010010110;
11'd1220 : tab = 23'b01000000110100000000100;
11'd1221 : tab = 23'b01000000101101101110101;
11'd1222 : tab = 23'b01000000100111011101000;
11'd1223 : tab = 23'b01000000100001001011100;
11'd1224 : tab = 23'b01000000011010111010011;
11'd1225 : tab = 23'b01000000010100101001011;
11'd1226 : tab = 23'b01000000001110011000110;
11'd1227 : tab = 23'b01000000001000001000010;
11'd1228 : tab = 23'b01000000000001111000001;
11'd1229 : tab = 23'b00111111111011101000001;
11'd1230 : tab = 23'b00111111110101011000100;
11'd1231 : tab = 23'b00111111101111001001000;
11'd1232 : tab = 23'b00111111101000111001110;
11'd1233 : tab = 23'b00111111100010101010110;
11'd1234 : tab = 23'b00111111011100011100000;
11'd1235 : tab = 23'b00111111010110001101100;
11'd1236 : tab = 23'b00111111001111111111010;
11'd1237 : tab = 23'b00111111001001110001010;
11'd1238 : tab = 23'b00111111000011100011100;
11'd1239 : tab = 23'b00111110111101010110000;
11'd1240 : tab = 23'b00111110110111001000110;
11'd1241 : tab = 23'b00111110110000111011110;
11'd1242 : tab = 23'b00111110101010101110111;
11'd1243 : tab = 23'b00111110100100100010010;
11'd1244 : tab = 23'b00111110011110010110000;
11'd1245 : tab = 23'b00111110011000001010000;
11'd1246 : tab = 23'b00111110010001111110000;
11'd1247 : tab = 23'b00111110001011110010100;
11'd1248 : tab = 23'b00111110000101100111010;
11'd1249 : tab = 23'b00111101111111011100000;
11'd1250 : tab = 23'b00111101111001010001010;
11'd1251 : tab = 23'b00111101110011000110100;
11'd1252 : tab = 23'b00111101101100111100001;
11'd1253 : tab = 23'b00111101100110110010000;
11'd1254 : tab = 23'b00111101100000101000000;
11'd1255 : tab = 23'b00111101011010011110011;
11'd1256 : tab = 23'b00111101010100010101000;
11'd1257 : tab = 23'b00111101001110001011110;
11'd1258 : tab = 23'b00111101001000000010110;
11'd1259 : tab = 23'b00111101000001111010000;
11'd1260 : tab = 23'b00111100111011110001100;
11'd1261 : tab = 23'b00111100110101101001010;
11'd1262 : tab = 23'b00111100101111100001010;
11'd1263 : tab = 23'b00111100101001011001100;
11'd1264 : tab = 23'b00111100100011010010000;
11'd1265 : tab = 23'b00111100011101001010110;
11'd1266 : tab = 23'b00111100010111000011100;
11'd1267 : tab = 23'b00111100010000111100110;
11'd1268 : tab = 23'b00111100001010110110010;
11'd1269 : tab = 23'b00111100000100101111110;
11'd1270 : tab = 23'b00111011111110101001110;
11'd1271 : tab = 23'b00111011111000100011110;
11'd1272 : tab = 23'b00111011110010011110001;
11'd1273 : tab = 23'b00111011101100011000110;
11'd1274 : tab = 23'b00111011100110010011100;
11'd1275 : tab = 23'b00111011100000001110100;
11'd1276 : tab = 23'b00111011011010001001111;
11'd1277 : tab = 23'b00111011010100000101011;
11'd1278 : tab = 23'b00111011001110000001001;
11'd1279 : tab = 23'b00111011000111111101000;
11'd1280 : tab = 23'b00111011000001111001010;
11'd1281 : tab = 23'b00111010111011110101110;
11'd1282 : tab = 23'b00111010110101110010100;
11'd1283 : tab = 23'b00111010101111101111010;
11'd1284 : tab = 23'b00111010101001101100100;
11'd1285 : tab = 23'b00111010100011101001110;
11'd1286 : tab = 23'b00111010011101100111100;
11'd1287 : tab = 23'b00111010010111100101010;
11'd1288 : tab = 23'b00111010010001100011011;
11'd1289 : tab = 23'b00111010001011100001101;
11'd1290 : tab = 23'b00111010000101100000010;
11'd1291 : tab = 23'b00111001111111011111000;
11'd1292 : tab = 23'b00111001111001011110000;
11'd1293 : tab = 23'b00111001110011011101010;
11'd1294 : tab = 23'b00111001101101011100101;
11'd1295 : tab = 23'b00111001100111011100010;
11'd1296 : tab = 23'b00111001100001011100010;
11'd1297 : tab = 23'b00111001011011011100011;
11'd1298 : tab = 23'b00111001010101011100110;
11'd1299 : tab = 23'b00111001001111011101011;
11'd1300 : tab = 23'b00111001001001011110010;
11'd1301 : tab = 23'b00111001000011011111010;
11'd1302 : tab = 23'b00111000111101100000100;
11'd1303 : tab = 23'b00111000110111100010000;
11'd1304 : tab = 23'b00111000110001100011110;
11'd1305 : tab = 23'b00111000101011100101110;
11'd1306 : tab = 23'b00111000100101101000000;
11'd1307 : tab = 23'b00111000011111101010100;
11'd1308 : tab = 23'b00111000011001101101000;
11'd1309 : tab = 23'b00111000010011110000000;
11'd1310 : tab = 23'b00111000001101110011000;
11'd1311 : tab = 23'b00111000000111110110011;
11'd1312 : tab = 23'b00111000000001111010000;
11'd1313 : tab = 23'b00110111111011111101110;
11'd1314 : tab = 23'b00110111110110000001110;
11'd1315 : tab = 23'b00110111110000000110000;
11'd1316 : tab = 23'b00110111101010001010100;
11'd1317 : tab = 23'b00110111100100001111010;
11'd1318 : tab = 23'b00110111011110010100000;
11'd1319 : tab = 23'b00110111011000011001010;
11'd1320 : tab = 23'b00110111010010011110101;
11'd1321 : tab = 23'b00110111001100100100010;
11'd1322 : tab = 23'b00110111000110101010000;
11'd1323 : tab = 23'b00110111000000110000000;
11'd1324 : tab = 23'b00110110111010110110011;
11'd1325 : tab = 23'b00110110110100111100110;
11'd1326 : tab = 23'b00110110101111000011100;
11'd1327 : tab = 23'b00110110101001001010100;
11'd1328 : tab = 23'b00110110100011010001110;
11'd1329 : tab = 23'b00110110011101011001000;
11'd1330 : tab = 23'b00110110010111100000101;
11'd1331 : tab = 23'b00110110010001101000100;
11'd1332 : tab = 23'b00110110001011110000100;
11'd1333 : tab = 23'b00110110000101111000110;
11'd1334 : tab = 23'b00110110000000000001010;
11'd1335 : tab = 23'b00110101111010001010000;
11'd1336 : tab = 23'b00110101110100010011000;
11'd1337 : tab = 23'b00110101101110011100000;
11'd1338 : tab = 23'b00110101101000100101100;
11'd1339 : tab = 23'b00110101100010101111001;
11'd1340 : tab = 23'b00110101011100111001000;
11'd1341 : tab = 23'b00110101010111000011000;
11'd1342 : tab = 23'b00110101010001001101010;
11'd1343 : tab = 23'b00110101001011010111110;
11'd1344 : tab = 23'b00110101000101100010100;
11'd1345 : tab = 23'b00110100111111101101010;
11'd1346 : tab = 23'b00110100111001111000100;
11'd1347 : tab = 23'b00110100110100000011111;
11'd1348 : tab = 23'b00110100101110001111100;
11'd1349 : tab = 23'b00110100101000011011010;
11'd1350 : tab = 23'b00110100100010100111010;
11'd1351 : tab = 23'b00110100011100110011100;
11'd1352 : tab = 23'b00110100010111000000000;
11'd1353 : tab = 23'b00110100010001001100110;
11'd1354 : tab = 23'b00110100001011011001100;
11'd1355 : tab = 23'b00110100000101100110110;
11'd1356 : tab = 23'b00110011111111110100000;
11'd1357 : tab = 23'b00110011111010000001101;
11'd1358 : tab = 23'b00110011110100001111011;
11'd1359 : tab = 23'b00110011101110011101011;
11'd1360 : tab = 23'b00110011101000101011100;
11'd1361 : tab = 23'b00110011100010111010000;
11'd1362 : tab = 23'b00110011011101001000101;
11'd1363 : tab = 23'b00110011010111010111100;
11'd1364 : tab = 23'b00110011010001100110100;
11'd1365 : tab = 23'b00110011001011110101111;
11'd1366 : tab = 23'b00110011000110000101011;
11'd1367 : tab = 23'b00110011000000010101000;
11'd1368 : tab = 23'b00110010111010100101000;
11'd1369 : tab = 23'b00110010110100110101010;
11'd1370 : tab = 23'b00110010101111000101100;
11'd1371 : tab = 23'b00110010101001010110001;
11'd1372 : tab = 23'b00110010100011100110111;
11'd1373 : tab = 23'b00110010011101110111111;
11'd1374 : tab = 23'b00110010011000001001001;
11'd1375 : tab = 23'b00110010010010011010100;
11'd1376 : tab = 23'b00110010001100101100010;
11'd1377 : tab = 23'b00110010000110111110000;
11'd1378 : tab = 23'b00110010000001010000001;
11'd1379 : tab = 23'b00110001111011100010100;
11'd1380 : tab = 23'b00110001110101110101000;
11'd1381 : tab = 23'b00110001110000000111110;
11'd1382 : tab = 23'b00110001101010011010100;
11'd1383 : tab = 23'b00110001100100101101110;
11'd1384 : tab = 23'b00110001011111000001001;
11'd1385 : tab = 23'b00110001011001010100110;
11'd1386 : tab = 23'b00110001010011101000100;
11'd1387 : tab = 23'b00110001001101111100100;
11'd1388 : tab = 23'b00110001001000010000110;
11'd1389 : tab = 23'b00110001000010100101000;
11'd1390 : tab = 23'b00110000111100111001110;
11'd1391 : tab = 23'b00110000110111001110100;
11'd1392 : tab = 23'b00110000110001100011101;
11'd1393 : tab = 23'b00110000101011111000111;
11'd1394 : tab = 23'b00110000100110001110011;
11'd1395 : tab = 23'b00110000100000100100000;
11'd1396 : tab = 23'b00110000011010111010000;
11'd1397 : tab = 23'b00110000010101010000000;
11'd1398 : tab = 23'b00110000001111100110011;
11'd1399 : tab = 23'b00110000001001111100111;
11'd1400 : tab = 23'b00110000000100010011101;
11'd1401 : tab = 23'b00101111111110101010100;
11'd1402 : tab = 23'b00101111111001000001110;
11'd1403 : tab = 23'b00101111110011011001001;
11'd1404 : tab = 23'b00101111101101110000101;
11'd1405 : tab = 23'b00101111101000001000100;
11'd1406 : tab = 23'b00101111100010100000100;
11'd1407 : tab = 23'b00101111011100111000110;
11'd1408 : tab = 23'b00101111010111010001000;
11'd1409 : tab = 23'b00101111010001101001101;
11'd1410 : tab = 23'b00101111001100000010100;
11'd1411 : tab = 23'b00101111000110011011100;
11'd1412 : tab = 23'b00101111000000110100110;
11'd1413 : tab = 23'b00101110111011001110010;
11'd1414 : tab = 23'b00101110110101100111110;
11'd1415 : tab = 23'b00101110110000000001110;
11'd1416 : tab = 23'b00101110101010011011110;
11'd1417 : tab = 23'b00101110100100110110000;
11'd1418 : tab = 23'b00101110011111010000100;
11'd1419 : tab = 23'b00101110011001101011010;
11'd1420 : tab = 23'b00101110010100000110000;
11'd1421 : tab = 23'b00101110001110100001010;
11'd1422 : tab = 23'b00101110001000111100100;
11'd1423 : tab = 23'b00101110000011011000000;
11'd1424 : tab = 23'b00101101111101110011110;
11'd1425 : tab = 23'b00101101111000001111101;
11'd1426 : tab = 23'b00101101110010101011110;
11'd1427 : tab = 23'b00101101101101001000000;
11'd1428 : tab = 23'b00101101100111100100101;
11'd1429 : tab = 23'b00101101100010000001010;
11'd1430 : tab = 23'b00101101011100011110010;
11'd1431 : tab = 23'b00101101010110111011100;
11'd1432 : tab = 23'b00101101010001011000110;
11'd1433 : tab = 23'b00101101001011110110011;
11'd1434 : tab = 23'b00101101000110010100000;
11'd1435 : tab = 23'b00101101000000110010000;
11'd1436 : tab = 23'b00101100111011010000010;
11'd1437 : tab = 23'b00101100110101101110100;
11'd1438 : tab = 23'b00101100110000001101001;
11'd1439 : tab = 23'b00101100101010101011111;
11'd1440 : tab = 23'b00101100100101001010111;
11'd1441 : tab = 23'b00101100011111101010000;
11'd1442 : tab = 23'b00101100011010001001100;
11'd1443 : tab = 23'b00101100010100101001000;
11'd1444 : tab = 23'b00101100001111001000110;
11'd1445 : tab = 23'b00101100001001101000110;
11'd1446 : tab = 23'b00101100000100001001000;
11'd1447 : tab = 23'b00101011111110101001011;
11'd1448 : tab = 23'b00101011111001001010000;
11'd1449 : tab = 23'b00101011110011101010110;
11'd1450 : tab = 23'b00101011101110001011110;
11'd1451 : tab = 23'b00101011101000101101000;
11'd1452 : tab = 23'b00101011100011001110010;
11'd1453 : tab = 23'b00101011011101101111111;
11'd1454 : tab = 23'b00101011011000010001110;
11'd1455 : tab = 23'b00101011010010110011110;
11'd1456 : tab = 23'b00101011001101010101110;
11'd1457 : tab = 23'b00101011000111111000010;
11'd1458 : tab = 23'b00101011000010011010111;
11'd1459 : tab = 23'b00101010111100111101101;
11'd1460 : tab = 23'b00101010110111100000101;
11'd1461 : tab = 23'b00101010110010000011110;
11'd1462 : tab = 23'b00101010101100100111010;
11'd1463 : tab = 23'b00101010100111001010110;
11'd1464 : tab = 23'b00101010100001101110100;
11'd1465 : tab = 23'b00101010011100010010100;
11'd1466 : tab = 23'b00101010010110110110110;
11'd1467 : tab = 23'b00101010010001011011001;
11'd1468 : tab = 23'b00101010001011111111101;
11'd1469 : tab = 23'b00101010000110100100100;
11'd1470 : tab = 23'b00101010000001001001100;
11'd1471 : tab = 23'b00101001111011101110100;
11'd1472 : tab = 23'b00101001110110010100000;
11'd1473 : tab = 23'b00101001110000111001100;
11'd1474 : tab = 23'b00101001101011011111010;
11'd1475 : tab = 23'b00101001100110000101010;
11'd1476 : tab = 23'b00101001100000101011011;
11'd1477 : tab = 23'b00101001011011010001110;
11'd1478 : tab = 23'b00101001010101111000010;
11'd1479 : tab = 23'b00101001010000011111000;
11'd1480 : tab = 23'b00101001001011000110000;
11'd1481 : tab = 23'b00101001000101101101000;
11'd1482 : tab = 23'b00101001000000010100011;
11'd1483 : tab = 23'b00101000111010111011111;
11'd1484 : tab = 23'b00101000110101100011100;
11'd1485 : tab = 23'b00101000110000001011100;
11'd1486 : tab = 23'b00101000101010110011101;
11'd1487 : tab = 23'b00101000100101011011111;
11'd1488 : tab = 23'b00101000100000000100100;
11'd1489 : tab = 23'b00101000011010101101000;
11'd1490 : tab = 23'b00101000010101010110000;
11'd1491 : tab = 23'b00101000001111111111000;
11'd1492 : tab = 23'b00101000001010101000010;
11'd1493 : tab = 23'b00101000000101010001110;
11'd1494 : tab = 23'b00100111111111111011100;
11'd1495 : tab = 23'b00100111111010100101010;
11'd1496 : tab = 23'b00100111110101001111011;
11'd1497 : tab = 23'b00100111101111111001100;
11'd1498 : tab = 23'b00100111101010100100000;
11'd1499 : tab = 23'b00100111100101001110101;
11'd1500 : tab = 23'b00100111011111111001011;
11'd1501 : tab = 23'b00100111011010100100100;
11'd1502 : tab = 23'b00100111010101001111110;
11'd1503 : tab = 23'b00100111001111111011000;
11'd1504 : tab = 23'b00100111001010100110101;
11'd1505 : tab = 23'b00100111000101010010011;
11'd1506 : tab = 23'b00100110111111111110010;
11'd1507 : tab = 23'b00100110111010101010100;
11'd1508 : tab = 23'b00100110110101010110111;
11'd1509 : tab = 23'b00100110110000000011011;
11'd1510 : tab = 23'b00100110101010110000000;
11'd1511 : tab = 23'b00100110100101011101000;
11'd1512 : tab = 23'b00100110100000001010001;
11'd1513 : tab = 23'b00100110011010110111100;
11'd1514 : tab = 23'b00100110010101100101000;
11'd1515 : tab = 23'b00100110010000010010100;
11'd1516 : tab = 23'b00100110001011000000100;
11'd1517 : tab = 23'b00100110000101101110100;
11'd1518 : tab = 23'b00100110000000011100110;
11'd1519 : tab = 23'b00100101111011001011010;
11'd1520 : tab = 23'b00100101110101111001111;
11'd1521 : tab = 23'b00100101110000101000101;
11'd1522 : tab = 23'b00100101101011010111110;
11'd1523 : tab = 23'b00100101100110000110110;
11'd1524 : tab = 23'b00100101100000110110010;
11'd1525 : tab = 23'b00100101011011100101110;
11'd1526 : tab = 23'b00100101010110010101100;
11'd1527 : tab = 23'b00100101010001000101100;
11'd1528 : tab = 23'b00100101001011110101101;
11'd1529 : tab = 23'b00100101000110100110000;
11'd1530 : tab = 23'b00100101000001010110100;
11'd1531 : tab = 23'b00100100111100000111010;
11'd1532 : tab = 23'b00100100110110111000000;
11'd1533 : tab = 23'b00100100110001101001001;
11'd1534 : tab = 23'b00100100101100011010011;
11'd1535 : tab = 23'b00100100100111001011110;
11'd1536 : tab = 23'b00100100100001111101100;
11'd1537 : tab = 23'b00100100011100101111010;
11'd1538 : tab = 23'b00100100010111100001010;
11'd1539 : tab = 23'b00100100010010010011100;
11'd1540 : tab = 23'b00100100001101000101111;
11'd1541 : tab = 23'b00100100000111111000100;
11'd1542 : tab = 23'b00100100000010101011010;
11'd1543 : tab = 23'b00100011111101011110001;
11'd1544 : tab = 23'b00100011111000010001010;
11'd1545 : tab = 23'b00100011110011000100100;
11'd1546 : tab = 23'b00100011101101111000000;
11'd1547 : tab = 23'b00100011101000101011110;
11'd1548 : tab = 23'b00100011100011011111100;
11'd1549 : tab = 23'b00100011011110010011101;
11'd1550 : tab = 23'b00100011011001000111110;
11'd1551 : tab = 23'b00100011010011111100010;
11'd1552 : tab = 23'b00100011001110110000111;
11'd1553 : tab = 23'b00100011001001100101101;
11'd1554 : tab = 23'b00100011000100011010100;
11'd1555 : tab = 23'b00100010111111001111110;
11'd1556 : tab = 23'b00100010111010000101001;
11'd1557 : tab = 23'b00100010110100111010101;
11'd1558 : tab = 23'b00100010101111110000010;
11'd1559 : tab = 23'b00100010101010100110010;
11'd1560 : tab = 23'b00100010100101011100010;
11'd1561 : tab = 23'b00100010100000010010100;
11'd1562 : tab = 23'b00100010011011001001000;
11'd1563 : tab = 23'b00100010010101111111100;
11'd1564 : tab = 23'b00100010010000110110011;
11'd1565 : tab = 23'b00100010001011101101010;
11'd1566 : tab = 23'b00100010000110100100100;
11'd1567 : tab = 23'b00100010000001011011111;
11'd1568 : tab = 23'b00100001111100010011011;
11'd1569 : tab = 23'b00100001110111001011000;
11'd1570 : tab = 23'b00100001110010000011000;
11'd1571 : tab = 23'b00100001101100111011000;
11'd1572 : tab = 23'b00100001100111110011010;
11'd1573 : tab = 23'b00100001100010101011110;
11'd1574 : tab = 23'b00100001011101100100010;
11'd1575 : tab = 23'b00100001011000011101001;
11'd1576 : tab = 23'b00100001010011010110000;
11'd1577 : tab = 23'b00100001001110001111010;
11'd1578 : tab = 23'b00100001001001001000100;
11'd1579 : tab = 23'b00100001000100000010000;
11'd1580 : tab = 23'b00100000111110111011110;
11'd1581 : tab = 23'b00100000111001110101101;
11'd1582 : tab = 23'b00100000110100101111110;
11'd1583 : tab = 23'b00100000101111101010000;
11'd1584 : tab = 23'b00100000101010100100010;
11'd1585 : tab = 23'b00100000100101011110111;
11'd1586 : tab = 23'b00100000100000011001110;
11'd1587 : tab = 23'b00100000011011010100110;
11'd1588 : tab = 23'b00100000010110001111110;
11'd1589 : tab = 23'b00100000010001001011001;
11'd1590 : tab = 23'b00100000001100000110100;
11'd1591 : tab = 23'b00100000000111000010010;
11'd1592 : tab = 23'b00100000000001111110001;
11'd1593 : tab = 23'b00011111111100111010001;
11'd1594 : tab = 23'b00011111110111110110010;
11'd1595 : tab = 23'b00011111110010110010110;
11'd1596 : tab = 23'b00011111101101101111010;
11'd1597 : tab = 23'b00011111101000101100000;
11'd1598 : tab = 23'b00011111100011101000111;
11'd1599 : tab = 23'b00011111011110100110000;
11'd1600 : tab = 23'b00011111011001100011010;
11'd1601 : tab = 23'b00011111010100100000110;
11'd1602 : tab = 23'b00011111001111011110010;
11'd1603 : tab = 23'b00011111001010011100000;
11'd1604 : tab = 23'b00011111000101011010000;
11'd1605 : tab = 23'b00011111000000011000010;
11'd1606 : tab = 23'b00011110111011010110100;
11'd1607 : tab = 23'b00011110110110010101000;
11'd1608 : tab = 23'b00011110110001010011110;
11'd1609 : tab = 23'b00011110101100010010100;
11'd1610 : tab = 23'b00011110100111010001100;
11'd1611 : tab = 23'b00011110100010010000110;
11'd1612 : tab = 23'b00011110011101010000001;
11'd1613 : tab = 23'b00011110011000001111101;
11'd1614 : tab = 23'b00011110010011001111011;
11'd1615 : tab = 23'b00011110001110001111010;
11'd1616 : tab = 23'b00011110001001001111011;
11'd1617 : tab = 23'b00011110000100001111100;
11'd1618 : tab = 23'b00011101111111010000000;
11'd1619 : tab = 23'b00011101111010010000101;
11'd1620 : tab = 23'b00011101110101010001011;
11'd1621 : tab = 23'b00011101110000010010010;
11'd1622 : tab = 23'b00011101101011010011100;
11'd1623 : tab = 23'b00011101100110010100110;
11'd1624 : tab = 23'b00011101100001010110010;
11'd1625 : tab = 23'b00011101011100010111111;
11'd1626 : tab = 23'b00011101010111011001101;
11'd1627 : tab = 23'b00011101010010011011110;
11'd1628 : tab = 23'b00011101001101011101110;
11'd1629 : tab = 23'b00011101001000100000001;
11'd1630 : tab = 23'b00011101000011100010110;
11'd1631 : tab = 23'b00011100111110100101010;
11'd1632 : tab = 23'b00011100111001101000010;
11'd1633 : tab = 23'b00011100110100101011010;
11'd1634 : tab = 23'b00011100101111101110100;
11'd1635 : tab = 23'b00011100101010110001110;
11'd1636 : tab = 23'b00011100100101110101010;
11'd1637 : tab = 23'b00011100100000111001000;
11'd1638 : tab = 23'b00011100011011111100111;
11'd1639 : tab = 23'b00011100010111000001000;
11'd1640 : tab = 23'b00011100010010000101010;
11'd1641 : tab = 23'b00011100001101001001100;
11'd1642 : tab = 23'b00011100001000001110001;
11'd1643 : tab = 23'b00011100000011010010111;
11'd1644 : tab = 23'b00011011111110010111110;
11'd1645 : tab = 23'b00011011111001011100111;
11'd1646 : tab = 23'b00011011110100100010001;
11'd1647 : tab = 23'b00011011101111100111100;
11'd1648 : tab = 23'b00011011101010101101001;
11'd1649 : tab = 23'b00011011100101110010111;
11'd1650 : tab = 23'b00011011100000111000110;
11'd1651 : tab = 23'b00011011011011111110111;
11'd1652 : tab = 23'b00011011010111000101010;
11'd1653 : tab = 23'b00011011010010001011101;
11'd1654 : tab = 23'b00011011001101010010010;
11'd1655 : tab = 23'b00011011001000011001000;
11'd1656 : tab = 23'b00011011000011100000000;
11'd1657 : tab = 23'b00011010111110100111001;
11'd1658 : tab = 23'b00011010111001101110011;
11'd1659 : tab = 23'b00011010110100110101110;
11'd1660 : tab = 23'b00011010101111111101100;
11'd1661 : tab = 23'b00011010101011000101010;
11'd1662 : tab = 23'b00011010100110001101010;
11'd1663 : tab = 23'b00011010100001010101010;
11'd1664 : tab = 23'b00011010011100011101101;
11'd1665 : tab = 23'b00011010010111100110000;
11'd1666 : tab = 23'b00011010010010101110110;
11'd1667 : tab = 23'b00011010001101110111100;
11'd1668 : tab = 23'b00011010001001000000100;
11'd1669 : tab = 23'b00011010000100001001101;
11'd1670 : tab = 23'b00011001111111010010111;
11'd1671 : tab = 23'b00011001111010011100010;
11'd1672 : tab = 23'b00011001110101100110000;
11'd1673 : tab = 23'b00011001110000101111110;
11'd1674 : tab = 23'b00011001101011111001110;
11'd1675 : tab = 23'b00011001100111000011111;
11'd1676 : tab = 23'b00011001100010001110010;
11'd1677 : tab = 23'b00011001011101011000110;
11'd1678 : tab = 23'b00011001011000100011010;
11'd1679 : tab = 23'b00011001010011101110001;
11'd1680 : tab = 23'b00011001001110111001000;
11'd1681 : tab = 23'b00011001001010000100010;
11'd1682 : tab = 23'b00011001000101001111100;
11'd1683 : tab = 23'b00011001000000011011000;
11'd1684 : tab = 23'b00011000111011100110100;
11'd1685 : tab = 23'b00011000110110110010011;
11'd1686 : tab = 23'b00011000110001111110010;
11'd1687 : tab = 23'b00011000101101001010100;
11'd1688 : tab = 23'b00011000101000010110110;
11'd1689 : tab = 23'b00011000100011100011010;
11'd1690 : tab = 23'b00011000011110101111110;
11'd1691 : tab = 23'b00011000011001111100100;
11'd1692 : tab = 23'b00011000010101001001100;
11'd1693 : tab = 23'b00011000010000010110101;
11'd1694 : tab = 23'b00011000001011100100000;
11'd1695 : tab = 23'b00011000000110110001010;
11'd1696 : tab = 23'b00011000000001111111000;
11'd1697 : tab = 23'b00010111111101001100110;
11'd1698 : tab = 23'b00010111111000011010101;
11'd1699 : tab = 23'b00010111110011101000110;
11'd1700 : tab = 23'b00010111101110110111000;
11'd1701 : tab = 23'b00010111101010000101011;
11'd1702 : tab = 23'b00010111100101010100000;
11'd1703 : tab = 23'b00010111100000100010110;
11'd1704 : tab = 23'b00010111011011110001101;
11'd1705 : tab = 23'b00010111010111000000110;
11'd1706 : tab = 23'b00010111010010010000000;
11'd1707 : tab = 23'b00010111001101011111010;
11'd1708 : tab = 23'b00010111001000101110111;
11'd1709 : tab = 23'b00010111000011111110100;
11'd1710 : tab = 23'b00010110111111001110100;
11'd1711 : tab = 23'b00010110111010011110100;
11'd1712 : tab = 23'b00010110110101101110110;
11'd1713 : tab = 23'b00010110110000111111001;
11'd1714 : tab = 23'b00010110101100001111101;
11'd1715 : tab = 23'b00010110100111100000010;
11'd1716 : tab = 23'b00010110100010110001001;
11'd1717 : tab = 23'b00010110011110000010010;
11'd1718 : tab = 23'b00010110011001010011010;
11'd1719 : tab = 23'b00010110010100100100101;
11'd1720 : tab = 23'b00010110001111110110010;
11'd1721 : tab = 23'b00010110001011000111110;
11'd1722 : tab = 23'b00010110000110011001101;
11'd1723 : tab = 23'b00010110000001101011100;
11'd1724 : tab = 23'b00010101111100111101110;
11'd1725 : tab = 23'b00010101111000010000000;
11'd1726 : tab = 23'b00010101110011100010100;
11'd1727 : tab = 23'b00010101101110110101000;
11'd1728 : tab = 23'b00010101101010000111110;
11'd1729 : tab = 23'b00010101100101011010110;
11'd1730 : tab = 23'b00010101100000101101111;
11'd1731 : tab = 23'b00010101011100000001000;
11'd1732 : tab = 23'b00010101010111010100100;
11'd1733 : tab = 23'b00010101010010101000001;
11'd1734 : tab = 23'b00010101001101111011110;
11'd1735 : tab = 23'b00010101001001001111110;
11'd1736 : tab = 23'b00010101000100100011110;
11'd1737 : tab = 23'b00010100111111111000000;
11'd1738 : tab = 23'b00010100111011001100010;
11'd1739 : tab = 23'b00010100110110100000110;
11'd1740 : tab = 23'b00010100110001110101100;
11'd1741 : tab = 23'b00010100101101001010011;
11'd1742 : tab = 23'b00010100101000011111010;
11'd1743 : tab = 23'b00010100100011110100100;
11'd1744 : tab = 23'b00010100011111001001110;
11'd1745 : tab = 23'b00010100011010011111010;
11'd1746 : tab = 23'b00010100010101110100111;
11'd1747 : tab = 23'b00010100010001001010110;
11'd1748 : tab = 23'b00010100001100100000100;
11'd1749 : tab = 23'b00010100000111110110110;
11'd1750 : tab = 23'b00010100000011001101000;
11'd1751 : tab = 23'b00010011111110100011011;
11'd1752 : tab = 23'b00010011111001111001111;
11'd1753 : tab = 23'b00010011110101010000110;
11'd1754 : tab = 23'b00010011110000100111100;
11'd1755 : tab = 23'b00010011101011111110100;
11'd1756 : tab = 23'b00010011100111010101110;
11'd1757 : tab = 23'b00010011100010101101001;
11'd1758 : tab = 23'b00010011011110000100100;
11'd1759 : tab = 23'b00010011011001011100010;
11'd1760 : tab = 23'b00010011010100110100000;
11'd1761 : tab = 23'b00010011010000001100000;
11'd1762 : tab = 23'b00010011001011100100001;
11'd1763 : tab = 23'b00010011000110111100100;
11'd1764 : tab = 23'b00010011000010010100110;
11'd1765 : tab = 23'b00010010111101101101100;
11'd1766 : tab = 23'b00010010111001000110010;
11'd1767 : tab = 23'b00010010110100011111001;
11'd1768 : tab = 23'b00010010101111111000001;
11'd1769 : tab = 23'b00010010101011010001010;
11'd1770 : tab = 23'b00010010100110101010110;
11'd1771 : tab = 23'b00010010100010000100010;
11'd1772 : tab = 23'b00010010011101011101111;
11'd1773 : tab = 23'b00010010011000110111110;
11'd1774 : tab = 23'b00010010010100010001110;
11'd1775 : tab = 23'b00010010001111101011111;
11'd1776 : tab = 23'b00010010001011000110001;
11'd1777 : tab = 23'b00010010000110100000100;
11'd1778 : tab = 23'b00010010000001111011001;
11'd1779 : tab = 23'b00010001111101010110000;
11'd1780 : tab = 23'b00010001111000110000110;
11'd1781 : tab = 23'b00010001110100001011111;
11'd1782 : tab = 23'b00010001101111100111000;
11'd1783 : tab = 23'b00010001101011000010011;
11'd1784 : tab = 23'b00010001100110011110000;
11'd1785 : tab = 23'b00010001100001111001101;
11'd1786 : tab = 23'b00010001011101010101011;
11'd1787 : tab = 23'b00010001011000110001011;
11'd1788 : tab = 23'b00010001010100001101100;
11'd1789 : tab = 23'b00010001001111101001110;
11'd1790 : tab = 23'b00010001001011000110010;
11'd1791 : tab = 23'b00010001000110100010110;
11'd1792 : tab = 23'b00010001000001111111100;
11'd1793 : tab = 23'b00010000111101011100011;
11'd1794 : tab = 23'b00010000111000111001100;
11'd1795 : tab = 23'b00010000110100010110100;
11'd1796 : tab = 23'b00010000101111110100000;
11'd1797 : tab = 23'b00010000101011010001100;
11'd1798 : tab = 23'b00010000100110101111000;
11'd1799 : tab = 23'b00010000100010001100111;
11'd1800 : tab = 23'b00010000011101101010110;
11'd1801 : tab = 23'b00010000011001001000111;
11'd1802 : tab = 23'b00010000010100100111000;
11'd1803 : tab = 23'b00010000010000000101100;
11'd1804 : tab = 23'b00010000001011100100000;
11'd1805 : tab = 23'b00010000000111000010110;
11'd1806 : tab = 23'b00010000000010100001101;
11'd1807 : tab = 23'b00001111111110000000100;
11'd1808 : tab = 23'b00001111111001011111110;
11'd1809 : tab = 23'b00001111110100111111000;
11'd1810 : tab = 23'b00001111110000011110100;
11'd1811 : tab = 23'b00001111101011111110000;
11'd1812 : tab = 23'b00001111100111011101110;
11'd1813 : tab = 23'b00001111100010111101101;
11'd1814 : tab = 23'b00001111011110011101110;
11'd1815 : tab = 23'b00001111011001111101111;
11'd1816 : tab = 23'b00001111010101011110010;
11'd1817 : tab = 23'b00001111010000111110110;
11'd1818 : tab = 23'b00001111001100011111011;
11'd1819 : tab = 23'b00001111001000000000001;
11'd1820 : tab = 23'b00001111000011100001000;
11'd1821 : tab = 23'b00001110111111000010001;
11'd1822 : tab = 23'b00001110111010100011010;
11'd1823 : tab = 23'b00001110110110000100110;
11'd1824 : tab = 23'b00001110110001100110010;
11'd1825 : tab = 23'b00001110101101001000000;
11'd1826 : tab = 23'b00001110101000101001110;
11'd1827 : tab = 23'b00001110100100001011110;
11'd1828 : tab = 23'b00001110011111101101111;
11'd1829 : tab = 23'b00001110011011010000000;
11'd1830 : tab = 23'b00001110010110110010100;
11'd1831 : tab = 23'b00001110010010010101000;
11'd1832 : tab = 23'b00001110001101110111110;
11'd1833 : tab = 23'b00001110001001011010101;
11'd1834 : tab = 23'b00001110000100111101100;
11'd1835 : tab = 23'b00001110000000100000110;
11'd1836 : tab = 23'b00001101111100000100000;
11'd1837 : tab = 23'b00001101110111100111100;
11'd1838 : tab = 23'b00001101110011001011000;
11'd1839 : tab = 23'b00001101101110101110110;
11'd1840 : tab = 23'b00001101101010010010101;
11'd1841 : tab = 23'b00001101100101110110110;
11'd1842 : tab = 23'b00001101100001011010111;
11'd1843 : tab = 23'b00001101011100111111010;
11'd1844 : tab = 23'b00001101011000100011101;
11'd1845 : tab = 23'b00001101010100001000010;
11'd1846 : tab = 23'b00001101001111101101000;
11'd1847 : tab = 23'b00001101001011010001111;
11'd1848 : tab = 23'b00001101000110110111000;
11'd1849 : tab = 23'b00001101000010011100001;
11'd1850 : tab = 23'b00001100111110000001100;
11'd1851 : tab = 23'b00001100111001100111000;
11'd1852 : tab = 23'b00001100110101001100100;
11'd1853 : tab = 23'b00001100110000110010010;
11'd1854 : tab = 23'b00001100101100011000010;
11'd1855 : tab = 23'b00001100100111111110010;
11'd1856 : tab = 23'b00001100100011100100100;
11'd1857 : tab = 23'b00001100011111001010111;
11'd1858 : tab = 23'b00001100011010110001010;
11'd1859 : tab = 23'b00001100010110011000000;
11'd1860 : tab = 23'b00001100010001111110110;
11'd1861 : tab = 23'b00001100001101100101101;
11'd1862 : tab = 23'b00001100001001001100110;
11'd1863 : tab = 23'b00001100000100110100000;
11'd1864 : tab = 23'b00001100000000011011010;
11'd1865 : tab = 23'b00001011111100000010110;
11'd1866 : tab = 23'b00001011110111101010011;
11'd1867 : tab = 23'b00001011110011010010010;
11'd1868 : tab = 23'b00001011101110111010001;
11'd1869 : tab = 23'b00001011101010100010010;
11'd1870 : tab = 23'b00001011100110001010100;
11'd1871 : tab = 23'b00001011100001110010110;
11'd1872 : tab = 23'b00001011011101011011010;
11'd1873 : tab = 23'b00001011011001000011111;
11'd1874 : tab = 23'b00001011010100101100110;
11'd1875 : tab = 23'b00001011010000010101100;
11'd1876 : tab = 23'b00001011001011111110101;
11'd1877 : tab = 23'b00001011000111100111110;
11'd1878 : tab = 23'b00001011000011010001010;
11'd1879 : tab = 23'b00001010111110111010110;
11'd1880 : tab = 23'b00001010111010100100011;
11'd1881 : tab = 23'b00001010110110001110001;
11'd1882 : tab = 23'b00001010110001111000000;
11'd1883 : tab = 23'b00001010101101100010000;
11'd1884 : tab = 23'b00001010101001001100010;
11'd1885 : tab = 23'b00001010100100110110101;
11'd1886 : tab = 23'b00001010100000100001000;
11'd1887 : tab = 23'b00001010011100001011110;
11'd1888 : tab = 23'b00001010010111110110100;
11'd1889 : tab = 23'b00001010010011100001011;
11'd1890 : tab = 23'b00001010001111001100100;
11'd1891 : tab = 23'b00001010001010110111101;
11'd1892 : tab = 23'b00001010000110100011000;
11'd1893 : tab = 23'b00001010000010001110100;
11'd1894 : tab = 23'b00001001111101111010000;
11'd1895 : tab = 23'b00001001111001100101110;
11'd1896 : tab = 23'b00001001110101010001101;
11'd1897 : tab = 23'b00001001110000111101110;
11'd1898 : tab = 23'b00001001101100101001111;
11'd1899 : tab = 23'b00001001101000010110010;
11'd1900 : tab = 23'b00001001100100000010101;
11'd1901 : tab = 23'b00001001011111101111010;
11'd1902 : tab = 23'b00001001011011011100000;
11'd1903 : tab = 23'b00001001010111001000110;
11'd1904 : tab = 23'b00001001010010110101110;
11'd1905 : tab = 23'b00001001001110100011000;
11'd1906 : tab = 23'b00001001001010010000010;
11'd1907 : tab = 23'b00001001000101111101101;
11'd1908 : tab = 23'b00001001000001101011010;
11'd1909 : tab = 23'b00001000111101011001000;
11'd1910 : tab = 23'b00001000111001000110110;
11'd1911 : tab = 23'b00001000110100110100110;
11'd1912 : tab = 23'b00001000110000100010111;
11'd1913 : tab = 23'b00001000101100010001000;
11'd1914 : tab = 23'b00001000100111111111100;
11'd1915 : tab = 23'b00001000100011101110000;
11'd1916 : tab = 23'b00001000011111011100110;
11'd1917 : tab = 23'b00001000011011001011100;
11'd1918 : tab = 23'b00001000010110111010100;
11'd1919 : tab = 23'b00001000010010101001100;
11'd1920 : tab = 23'b00001000001110011000110;
11'd1921 : tab = 23'b00001000001010001000000;
11'd1922 : tab = 23'b00001000000101110111100;
11'd1923 : tab = 23'b00001000000001100111010;
11'd1924 : tab = 23'b00000111111101010111000;
11'd1925 : tab = 23'b00000111111001000110111;
11'd1926 : tab = 23'b00000111110100110110111;
11'd1927 : tab = 23'b00000111110000100111000;
11'd1928 : tab = 23'b00000111101100010111011;
11'd1929 : tab = 23'b00000111101000000111110;
11'd1930 : tab = 23'b00000111100011111000100;
11'd1931 : tab = 23'b00000111011111101001010;
11'd1932 : tab = 23'b00000111011011011010000;
11'd1933 : tab = 23'b00000111010111001011000;
11'd1934 : tab = 23'b00000111010010111100001;
11'd1935 : tab = 23'b00000111001110101101100;
11'd1936 : tab = 23'b00000111001010011110110;
11'd1937 : tab = 23'b00000111000110010000010;
11'd1938 : tab = 23'b00000111000010000010000;
11'd1939 : tab = 23'b00000110111101110011110;
11'd1940 : tab = 23'b00000110111001100101110;
11'd1941 : tab = 23'b00000110110101010111111;
11'd1942 : tab = 23'b00000110110001001010000;
11'd1943 : tab = 23'b00000110101100111100100;
11'd1944 : tab = 23'b00000110101000101111000;
11'd1945 : tab = 23'b00000110100100100001100;
11'd1946 : tab = 23'b00000110100000010100010;
11'd1947 : tab = 23'b00000110011100000111010;
11'd1948 : tab = 23'b00000110010111111010010;
11'd1949 : tab = 23'b00000110010011101101011;
11'd1950 : tab = 23'b00000110001111100000110;
11'd1951 : tab = 23'b00000110001011010100001;
11'd1952 : tab = 23'b00000110000111000111110;
11'd1953 : tab = 23'b00000110000010111011011;
11'd1954 : tab = 23'b00000101111110101111010;
11'd1955 : tab = 23'b00000101111010100011010;
11'd1956 : tab = 23'b00000101110110010111010;
11'd1957 : tab = 23'b00000101110010001011100;
11'd1958 : tab = 23'b00000101101101111111111;
11'd1959 : tab = 23'b00000101101001110100011;
11'd1960 : tab = 23'b00000101100101101001000;
11'd1961 : tab = 23'b00000101100001011101110;
11'd1962 : tab = 23'b00000101011101010010110;
11'd1963 : tab = 23'b00000101011001000111110;
11'd1964 : tab = 23'b00000101010100111100111;
11'd1965 : tab = 23'b00000101010000110010010;
11'd1966 : tab = 23'b00000101001100100111101;
11'd1967 : tab = 23'b00000101001000011101010;
11'd1968 : tab = 23'b00000101000100010010111;
11'd1969 : tab = 23'b00000101000000001000110;
11'd1970 : tab = 23'b00000100111011111110110;
11'd1971 : tab = 23'b00000100110111110100110;
11'd1972 : tab = 23'b00000100110011101011000;
11'd1973 : tab = 23'b00000100101111100001011;
11'd1974 : tab = 23'b00000100101011010111110;
11'd1975 : tab = 23'b00000100100111001110100;
11'd1976 : tab = 23'b00000100100011000101010;
11'd1977 : tab = 23'b00000100011110111100001;
11'd1978 : tab = 23'b00000100011010110011010;
11'd1979 : tab = 23'b00000100010110101010010;
11'd1980 : tab = 23'b00000100010010100001100;
11'd1981 : tab = 23'b00000100001110011001000;
11'd1982 : tab = 23'b00000100001010010000100;
11'd1983 : tab = 23'b00000100000110001000010;
11'd1984 : tab = 23'b00000100000010000000000;
11'd1985 : tab = 23'b00000011111101111000000;
11'd1986 : tab = 23'b00000011111001110000000;
11'd1987 : tab = 23'b00000011110101101000010;
11'd1988 : tab = 23'b00000011110001100000100;
11'd1989 : tab = 23'b00000011101101011001000;
11'd1990 : tab = 23'b00000011101001010001101;
11'd1991 : tab = 23'b00000011100101001010010;
11'd1992 : tab = 23'b00000011100001000011010;
11'd1993 : tab = 23'b00000011011100111100010;
11'd1994 : tab = 23'b00000011011000110101010;
11'd1995 : tab = 23'b00000011010100101110100;
11'd1996 : tab = 23'b00000011010000100111111;
11'd1997 : tab = 23'b00000011001100100001100;
11'd1998 : tab = 23'b00000011001000011011000;
11'd1999 : tab = 23'b00000011000100010100110;
11'd2000 : tab = 23'b00000011000000001110110;
11'd2001 : tab = 23'b00000010111100001000110;
11'd2002 : tab = 23'b00000010111000000010111;
11'd2003 : tab = 23'b00000010110011111101010;
11'd2004 : tab = 23'b00000010101111110111101;
11'd2005 : tab = 23'b00000010101011110010001;
11'd2006 : tab = 23'b00000010100111101100110;
11'd2007 : tab = 23'b00000010100011100111100;
11'd2008 : tab = 23'b00000010011111100010100;
11'd2009 : tab = 23'b00000010011011011101100;
11'd2010 : tab = 23'b00000010010111011000110;
11'd2011 : tab = 23'b00000010010011010100000;
11'd2012 : tab = 23'b00000010001111001111100;
11'd2013 : tab = 23'b00000010001011001011000;
11'd2014 : tab = 23'b00000010000111000110110;
11'd2015 : tab = 23'b00000010000011000010101;
11'd2016 : tab = 23'b00000001111110111110100;
11'd2017 : tab = 23'b00000001111010111010101;
11'd2018 : tab = 23'b00000001110110110110110;
11'd2019 : tab = 23'b00000001110010110011001;
11'd2020 : tab = 23'b00000001101110101111101;
11'd2021 : tab = 23'b00000001101010101100010;
11'd2022 : tab = 23'b00000001100110101001000;
11'd2023 : tab = 23'b00000001100010100101110;
11'd2024 : tab = 23'b00000001011110100010110;
11'd2025 : tab = 23'b00000001011010011111111;
11'd2026 : tab = 23'b00000001010110011101000;
11'd2027 : tab = 23'b00000001010010011010100;
11'd2028 : tab = 23'b00000001001110011000000;
11'd2029 : tab = 23'b00000001001010010101100;
11'd2030 : tab = 23'b00000001000110010011010;
11'd2031 : tab = 23'b00000001000010010001001;
11'd2032 : tab = 23'b00000000111110001111001;
11'd2033 : tab = 23'b00000000111010001101010;
11'd2034 : tab = 23'b00000000110110001011100;
11'd2035 : tab = 23'b00000000110010001001111;
11'd2036 : tab = 23'b00000000101110001000010;
11'd2037 : tab = 23'b00000000101010000111000;
11'd2038 : tab = 23'b00000000100110000101110;
11'd2039 : tab = 23'b00000000100010000100101;
11'd2040 : tab = 23'b00000000011110000011100;
11'd2041 : tab = 23'b00000000011010000010110;
11'd2042 : tab = 23'b00000000010110000010000;
11'd2043 : tab = 23'b00000000010010000001011;
11'd2044 : tab = 23'b00000000001110000000110;
11'd2045 : tab = 23'b00000000001010000000100;
11'd2046 : tab = 23'b00000000000110000000010;
11'd2047 : tab = 23'b00000000000010000000001;
endcase
  end
  endfunction
  
  function [22:0] tab2 (
    input [10:0] N
  );
  begin
  case(N)
11'd0 : tab2 = 23'b11111111110000000000111;
11'd1 : tab2 = 23'b11111111010000000011111;
11'd2 : tab2 = 23'b11111110110000001001111;
11'd3 : tab2 = 23'b11111110010000010010111;
11'd4 : tab2 = 23'b11111101110000011110111;
11'd5 : tab2 = 23'b11111101010000101101110;
11'd6 : tab2 = 23'b11111100110000111111100;
11'd7 : tab2 = 23'b11111100010001010100011;
11'd8 : tab2 = 23'b11111011110001101100011;
11'd9 : tab2 = 23'b11111011010010000111010;
11'd10 : tab2 = 23'b11111010110010100100100;
11'd11 : tab2 = 23'b11111010010011000101011;
11'd12 : tab2 = 23'b11111001110011101001001;
11'd13 : tab2 = 23'b11111001010100001111011;
11'd14 : tab2 = 23'b11111000110100111000111;
11'd15 : tab2 = 23'b11111000010101100101011;
11'd16 : tab2 = 23'b11110111110110010100100;
11'd17 : tab2 = 23'b11110111010111000110100;
11'd18 : tab2 = 23'b11110110110111111011111;
11'd19 : tab2 = 23'b11110110011000110011100;
11'd20 : tab2 = 23'b11110101111001101110100;
11'd21 : tab2 = 23'b11110101011010101100011;
11'd22 : tab2 = 23'b11110100111011101100101;
11'd23 : tab2 = 23'b11110100011100110000011;
11'd24 : tab2 = 23'b11110011111101110110101;
11'd25 : tab2 = 23'b11110011011110111111111;
11'd26 : tab2 = 23'b11110011000000001100000;
11'd27 : tab2 = 23'b11110010100001011010111;
11'd28 : tab2 = 23'b11110010000010101100100;
11'd29 : tab2 = 23'b11110001100100000001011;
11'd30 : tab2 = 23'b11110001000101011000101;
11'd31 : tab2 = 23'b11110000100110110011000;
11'd32 : tab2 = 23'b11110000001000010000000;
11'd33 : tab2 = 23'b11101111101001101111110;
11'd34 : tab2 = 23'b11101111001011010010100;
11'd35 : tab2 = 23'b11101110101100111000001;
11'd36 : tab2 = 23'b11101110001110100000100;
11'd37 : tab2 = 23'b11101101110000001011100;
11'd38 : tab2 = 23'b11101101010001111001100;
11'd39 : tab2 = 23'b11101100110011101001111;
11'd40 : tab2 = 23'b11101100010101011101101;
11'd41 : tab2 = 23'b11101011110111010011110;
11'd42 : tab2 = 23'b11101011011001001100110;
11'd43 : tab2 = 23'b11101010111011001000101;
11'd44 : tab2 = 23'b11101010011101000111000;
11'd45 : tab2 = 23'b11101001111111001000011;
11'd46 : tab2 = 23'b11101001100001001100011;
11'd47 : tab2 = 23'b11101001000011010011000;
11'd48 : tab2 = 23'b11101000100101011100101;
11'd49 : tab2 = 23'b11101000000111101001000;
11'd50 : tab2 = 23'b11100111101001111000000;
11'd51 : tab2 = 23'b11100111001100001001011;
11'd52 : tab2 = 23'b11100110101110011101111;
11'd53 : tab2 = 23'b11100110010000110101001;
11'd54 : tab2 = 23'b11100101110011001110101;
11'd55 : tab2 = 23'b11100101010101101011011;
11'd56 : tab2 = 23'b11100100111000001010100;
11'd57 : tab2 = 23'b11100100011010101100100;
11'd58 : tab2 = 23'b11100011111101010000111;
11'd59 : tab2 = 23'b11100011011111111000011;
11'd60 : tab2 = 23'b11100011000010100010001;
11'd61 : tab2 = 23'b11100010100101001111000;
11'd62 : tab2 = 23'b11100010000111111110001;
11'd63 : tab2 = 23'b11100001101010110000001;
11'd64 : tab2 = 23'b11100001001101100100110;
11'd65 : tab2 = 23'b11100000110000011100000;
11'd66 : tab2 = 23'b11100000010011010101110;
11'd67 : tab2 = 23'b11011111110110010010010;
11'd68 : tab2 = 23'b11011111011001010001110;
11'd69 : tab2 = 23'b11011110111100010011001;
11'd70 : tab2 = 23'b11011110011111010111110;
11'd71 : tab2 = 23'b11011110000010011110110;
11'd72 : tab2 = 23'b11011101100101101000100;
11'd73 : tab2 = 23'b11011101001000110100110;
11'd74 : tab2 = 23'b11011100101100000011110;
11'd75 : tab2 = 23'b11011100001111010101000;
11'd76 : tab2 = 23'b11011011110010101001001;
11'd77 : tab2 = 23'b11011011010101111111111;
11'd78 : tab2 = 23'b11011010111001011001001;
11'd79 : tab2 = 23'b11011010011100110100111;
11'd80 : tab2 = 23'b11011010000000010011001;
11'd81 : tab2 = 23'b11011001100011110100010;
11'd82 : tab2 = 23'b11011001000111010111111;
11'd83 : tab2 = 23'b11011000101010111101111;
11'd84 : tab2 = 23'b11011000001110100110100;
11'd85 : tab2 = 23'b11010111110010010001110;
11'd86 : tab2 = 23'b11010111010101111111100;
11'd87 : tab2 = 23'b11010110111001101111111;
11'd88 : tab2 = 23'b11010110011101100010101;
11'd89 : tab2 = 23'b11010110000001011000000;
11'd90 : tab2 = 23'b11010101100101001111111;
11'd91 : tab2 = 23'b11010101001001001010010;
11'd92 : tab2 = 23'b11010100101101000111011;
11'd93 : tab2 = 23'b11010100010001000110110;
11'd94 : tab2 = 23'b11010011110101001000101;
11'd95 : tab2 = 23'b11010011011001001101011;
11'd96 : tab2 = 23'b11010010111101010100000;
11'd97 : tab2 = 23'b11010010100001011101101;
11'd98 : tab2 = 23'b11010010000101101001101;
11'd99 : tab2 = 23'b11010001101001111000000;
11'd100 : tab2 = 23'b11010001001110001001000;
11'd101 : tab2 = 23'b11010000110010011100001;
11'd102 : tab2 = 23'b11010000010110110010010;
11'd103 : tab2 = 23'b11001111111011001010101;
11'd104 : tab2 = 23'b11001111011111100101011;
11'd105 : tab2 = 23'b11001111000100000010101;
11'd106 : tab2 = 23'b11001110101000100010010;
11'd107 : tab2 = 23'b11001110001101000100101;
11'd108 : tab2 = 23'b11001101110001101001010;
11'd109 : tab2 = 23'b11001101010110010000000;
11'd110 : tab2 = 23'b11001100111010111001100;
11'd111 : tab2 = 23'b11001100011111100101100;
11'd112 : tab2 = 23'b11001100000100010011110;
11'd113 : tab2 = 23'b11001011101001000100101;
11'd114 : tab2 = 23'b11001011001101110111111;
11'd115 : tab2 = 23'b11001010110010101101011;
11'd116 : tab2 = 23'b11001010010111100101100;
11'd117 : tab2 = 23'b11001001111100011111110;
11'd118 : tab2 = 23'b11001001100001011100100;
11'd119 : tab2 = 23'b11001001000110011100000;
11'd120 : tab2 = 23'b11001000101011011101101;
11'd121 : tab2 = 23'b11001000010000100001100;
11'd122 : tab2 = 23'b11000111110101100111111;
11'd123 : tab2 = 23'b11000111011010110000101;
11'd124 : tab2 = 23'b11000110111111111011110;
11'd125 : tab2 = 23'b11000110100101001001001;
11'd126 : tab2 = 23'b11000110001010011001000;
11'd127 : tab2 = 23'b11000101101111101011010;
11'd128 : tab2 = 23'b11000101010100111111110;
11'd129 : tab2 = 23'b11000100111010010110111;
11'd130 : tab2 = 23'b11000100011111110000000;
11'd131 : tab2 = 23'b11000100000101001011110;
11'd132 : tab2 = 23'b11000011101010101001101;
11'd133 : tab2 = 23'b11000011010000001001111;
11'd134 : tab2 = 23'b11000010110101101100101;
11'd135 : tab2 = 23'b11000010011011010001101;
11'd136 : tab2 = 23'b11000010000000111000110;
11'd137 : tab2 = 23'b11000001100110100010010;
11'd138 : tab2 = 23'b11000001001100001110000;
11'd139 : tab2 = 23'b11000000110001111100001;
11'd140 : tab2 = 23'b11000000010111101101000;
11'd141 : tab2 = 23'b10111111111101011111101;
11'd142 : tab2 = 23'b10111111100011010100101;
11'd143 : tab2 = 23'b10111111001001001100001;
11'd144 : tab2 = 23'b10111110101111000101110;
11'd145 : tab2 = 23'b10111110010101000001111;
11'd146 : tab2 = 23'b10111101111011000000001;
11'd147 : tab2 = 23'b10111101100001000000100;
11'd148 : tab2 = 23'b10111101000111000011011;
11'd149 : tab2 = 23'b10111100101101001000010;
11'd150 : tab2 = 23'b10111100010011001111101;
11'd151 : tab2 = 23'b10111011111001011001011;
11'd152 : tab2 = 23'b10111011011111100101010;
11'd153 : tab2 = 23'b10111011000101110011010;
11'd154 : tab2 = 23'b10111010101100000011101;
11'd155 : tab2 = 23'b10111010010010010110011;
11'd156 : tab2 = 23'b10111001111000101011001;
11'd157 : tab2 = 23'b10111001011111000010001;
11'd158 : tab2 = 23'b10111001000101011011010;
11'd159 : tab2 = 23'b10111000101011110110111;
11'd160 : tab2 = 23'b10111000010010010100100;
11'd161 : tab2 = 23'b10110111111000110100101;
11'd162 : tab2 = 23'b10110111011111010110110;
11'd163 : tab2 = 23'b10110111000101111011000;
11'd164 : tab2 = 23'b10110110101100100001110;
11'd165 : tab2 = 23'b10110110010011001010010;
11'd166 : tab2 = 23'b10110101111001110101101;
11'd167 : tab2 = 23'b10110101100000100010101;
11'd168 : tab2 = 23'b10110101000111010010000;
11'd169 : tab2 = 23'b10110100101110000011100;
11'd170 : tab2 = 23'b10110100010100110111010;
11'd171 : tab2 = 23'b10110011111011101101010;
11'd172 : tab2 = 23'b10110011100010100101010;
11'd173 : tab2 = 23'b10110011001001011111011;
11'd174 : tab2 = 23'b10110010110000011100001;
11'd175 : tab2 = 23'b10110010010111011010100;
11'd176 : tab2 = 23'b10110001111110011011011;
11'd177 : tab2 = 23'b10110001100101011110010;
11'd178 : tab2 = 23'b10110001001100100011011;
11'd179 : tab2 = 23'b10110000110011101010100;
11'd180 : tab2 = 23'b10110000011010110100001;
11'd181 : tab2 = 23'b10110000000001111111100;
11'd182 : tab2 = 23'b10101111101001001101000;
11'd183 : tab2 = 23'b10101111010000011100110;
11'd184 : tab2 = 23'b10101110110111101110101;
11'd185 : tab2 = 23'b10101110011111000010101;
11'd186 : tab2 = 23'b10101110000110011000110;
11'd187 : tab2 = 23'b10101101101101110001000;
11'd188 : tab2 = 23'b10101101010101001011100;
11'd189 : tab2 = 23'b10101100111100101000000;
11'd190 : tab2 = 23'b10101100100100000110011;
11'd191 : tab2 = 23'b10101100001011100111010;
11'd192 : tab2 = 23'b10101011110011001010000;
11'd193 : tab2 = 23'b10101011011010101110111;
11'd194 : tab2 = 23'b10101011000010010101110;
11'd195 : tab2 = 23'b10101010101001111110101;
11'd196 : tab2 = 23'b10101010010001101001111;
11'd197 : tab2 = 23'b10101001111001010111010;
11'd198 : tab2 = 23'b10101001100001000110011;
11'd199 : tab2 = 23'b10101001001000110111110;
11'd200 : tab2 = 23'b10101000110000101011010;
11'd201 : tab2 = 23'b10101000011000100000100;
11'd202 : tab2 = 23'b10101000000000011000011;
11'd203 : tab2 = 23'b10100111101000010001110;
11'd204 : tab2 = 23'b10100111010000001101101;
11'd205 : tab2 = 23'b10100110111000001011001;
11'd206 : tab2 = 23'b10100110100000001011001;
11'd207 : tab2 = 23'b10100110001000001100110;
11'd208 : tab2 = 23'b10100101110000010000101;
11'd209 : tab2 = 23'b10100101011000010110100;
11'd210 : tab2 = 23'b10100101000000011110011;
11'd211 : tab2 = 23'b10100100101000101000011;
11'd212 : tab2 = 23'b10100100010000110100001;
11'd213 : tab2 = 23'b10100011111001000010100;
11'd214 : tab2 = 23'b10100011100001010010010;
11'd215 : tab2 = 23'b10100011001001100100011;
11'd216 : tab2 = 23'b10100010110001111000100;
11'd217 : tab2 = 23'b10100010011010001110100;
11'd218 : tab2 = 23'b10100010000010100110011;
11'd219 : tab2 = 23'b10100001101011000000011;
11'd220 : tab2 = 23'b10100001010011011100011;
11'd221 : tab2 = 23'b10100000111011111010101;
11'd222 : tab2 = 23'b10100000100100011010101;
11'd223 : tab2 = 23'b10100000001100111100101;
11'd224 : tab2 = 23'b10011111110101100000100;
11'd225 : tab2 = 23'b10011111011110000110101;
11'd226 : tab2 = 23'b10011111000110101110011;
11'd227 : tab2 = 23'b10011110101111011000010;
11'd228 : tab2 = 23'b10011110011000000100011;
11'd229 : tab2 = 23'b10011110000000110010000;
11'd230 : tab2 = 23'b10011101101001100010001;
11'd231 : tab2 = 23'b10011101010010010011110;
11'd232 : tab2 = 23'b10011100111011000111011;
11'd233 : tab2 = 23'b10011100100011111101000;
11'd234 : tab2 = 23'b10011100001100110100110;
11'd235 : tab2 = 23'b10011011110101101110011;
11'd236 : tab2 = 23'b10011011011110101001110;
11'd237 : tab2 = 23'b10011011000111100111001;
11'd238 : tab2 = 23'b10011010110000100110110;
11'd239 : tab2 = 23'b10011010011001100111111;
11'd240 : tab2 = 23'b10011010000010101011000;
11'd241 : tab2 = 23'b10011001101011110000011;
11'd242 : tab2 = 23'b10011001010100110111100;
11'd243 : tab2 = 23'b10011000111110000000011;
11'd244 : tab2 = 23'b10011000100111001011011;
11'd245 : tab2 = 23'b10011000010000011000010;
11'd246 : tab2 = 23'b10010111111001100111000;
11'd247 : tab2 = 23'b10010111100010110111100;
11'd248 : tab2 = 23'b10010111001100001010000;
11'd249 : tab2 = 23'b10010110110101011110100;
11'd250 : tab2 = 23'b10010110011110110100110;
11'd251 : tab2 = 23'b10010110001000001100111;
11'd252 : tab2 = 23'b10010101110001100111010;
11'd253 : tab2 = 23'b10010101011011000011010;
11'd254 : tab2 = 23'b10010101000100100001000;
11'd255 : tab2 = 23'b10010100101110000000101;
11'd256 : tab2 = 23'b10010100010111100010011;
11'd257 : tab2 = 23'b10010100000001000101111;
11'd258 : tab2 = 23'b10010011101010101011001;
11'd259 : tab2 = 23'b10010011010100010010011;
11'd260 : tab2 = 23'b10010010111101111011100;
11'd261 : tab2 = 23'b10010010100111100110101;
11'd262 : tab2 = 23'b10010010010001010011010;
11'd263 : tab2 = 23'b10010001111011000001110;
11'd264 : tab2 = 23'b10010001100100110010100;
11'd265 : tab2 = 23'b10010001001110100100110;
11'd266 : tab2 = 23'b10010000111000011001001;
11'd267 : tab2 = 23'b10010000100010001111000;
11'd268 : tab2 = 23'b10010000001100000110111;
11'd269 : tab2 = 23'b10001111110110000000101;
11'd270 : tab2 = 23'b10001111011111111100010;
11'd271 : tab2 = 23'b10001111001001111001100;
11'd272 : tab2 = 23'b10001110110011111000101;
11'd273 : tab2 = 23'b10001110011101111001101;
11'd274 : tab2 = 23'b10001110000111111100101;
11'd275 : tab2 = 23'b10001101110010000001000;
11'd276 : tab2 = 23'b10001101011100000111100;
11'd277 : tab2 = 23'b10001101000110001111110;
11'd278 : tab2 = 23'b10001100110000011010000;
11'd279 : tab2 = 23'b10001100011010100101110;
11'd280 : tab2 = 23'b10001100000100110011011;
11'd281 : tab2 = 23'b10001011101111000010111;
11'd282 : tab2 = 23'b10001011011001010011111;
11'd283 : tab2 = 23'b10001011000011100111001;
11'd284 : tab2 = 23'b10001010101101111100000;
11'd285 : tab2 = 23'b10001010011000010010100;
11'd286 : tab2 = 23'b10001010000010101010110;
11'd287 : tab2 = 23'b10001001101101000100111;
11'd288 : tab2 = 23'b10001001010111100001000;
11'd289 : tab2 = 23'b10001001000001111110100;
11'd290 : tab2 = 23'b10001000101100011110001;
11'd291 : tab2 = 23'b10001000010110111111010;
11'd292 : tab2 = 23'b10001000000001100010100;
11'd293 : tab2 = 23'b10000111101100000111001;
11'd294 : tab2 = 23'b10000111010110101101100;
11'd295 : tab2 = 23'b10000111000001010101110;
11'd296 : tab2 = 23'b10000110101011111111110;
11'd297 : tab2 = 23'b10000110010110101011100;
11'd298 : tab2 = 23'b10000110000001011001010;
11'd299 : tab2 = 23'b10000101101100001000011;
11'd300 : tab2 = 23'b10000101010110111001010;
11'd301 : tab2 = 23'b10000101000001101100000;
11'd302 : tab2 = 23'b10000100101100100000011;
11'd303 : tab2 = 23'b10000100010111010110101;
11'd304 : tab2 = 23'b10000100000010001110011;
11'd305 : tab2 = 23'b10000011101101001000010;
11'd306 : tab2 = 23'b10000011011000000011100;
11'd307 : tab2 = 23'b10000011000011000000011;
11'd308 : tab2 = 23'b10000010101101111111100;
11'd309 : tab2 = 23'b10000010011000111111111;
11'd310 : tab2 = 23'b10000010000100000010000;
11'd311 : tab2 = 23'b10000001101111000110000;
11'd312 : tab2 = 23'b10000001011010001011100;
11'd313 : tab2 = 23'b10000001000101010011000;
11'd314 : tab2 = 23'b10000000110000011011111;
11'd315 : tab2 = 23'b10000000011011100110100;
11'd316 : tab2 = 23'b10000000000110110010111;
11'd317 : tab2 = 23'b01111111110010000001010;
11'd318 : tab2 = 23'b01111111011101010000110;
11'd319 : tab2 = 23'b01111111001000100010001;
11'd320 : tab2 = 23'b01111110110011110101011;
11'd321 : tab2 = 23'b01111110011111001010001;
11'd322 : tab2 = 23'b01111110001010100000110;
11'd323 : tab2 = 23'b01111101110101111000110;
11'd324 : tab2 = 23'b01111101100001010010100;
11'd325 : tab2 = 23'b01111101001100101110000;
11'd326 : tab2 = 23'b01111100111000001011010;
11'd327 : tab2 = 23'b01111100100011101010000;
11'd328 : tab2 = 23'b01111100001111001010100;
11'd329 : tab2 = 23'b01111011111010101100101;
11'd330 : tab2 = 23'b01111011100110010000100;
11'd331 : tab2 = 23'b01111011010001110101111;
11'd332 : tab2 = 23'b01111010111101011100111;
11'd333 : tab2 = 23'b01111010101001000101101;
11'd334 : tab2 = 23'b01111010010100110000001;
11'd335 : tab2 = 23'b01111010000000011011110;
11'd336 : tab2 = 23'b01111001101100001001100;
11'd337 : tab2 = 23'b01111001010111111000101;
11'd338 : tab2 = 23'b01111001000011101001101;
11'd339 : tab2 = 23'b01111000101111011100010;
11'd340 : tab2 = 23'b01111000011011010000100;
11'd341 : tab2 = 23'b01111000000111000110000;
11'd342 : tab2 = 23'b01110111110010111101100;
11'd343 : tab2 = 23'b01110111011110110110100;
11'd344 : tab2 = 23'b01110111001010110001000;
11'd345 : tab2 = 23'b01110110110110101101010;
11'd346 : tab2 = 23'b01110110100010101011010;
11'd347 : tab2 = 23'b01110110001110101010100;
11'd348 : tab2 = 23'b01110101111010101011101;
11'd349 : tab2 = 23'b01110101100110101110010;
11'd350 : tab2 = 23'b01110101010010110010011;
11'd351 : tab2 = 23'b01110100111110111000010;
11'd352 : tab2 = 23'b01110100101010111111101;
11'd353 : tab2 = 23'b01110100010111001000110;
11'd354 : tab2 = 23'b01110100000011010011011;
11'd355 : tab2 = 23'b01110011101111011111011;
11'd356 : tab2 = 23'b01110011011011101101010;
11'd357 : tab2 = 23'b01110011000111111100110;
11'd358 : tab2 = 23'b01110010110100001101100;
11'd359 : tab2 = 23'b01110010100000011111111;
11'd360 : tab2 = 23'b01110010001100110100001;
11'd361 : tab2 = 23'b01110001111001001001100;
11'd362 : tab2 = 23'b01110001100101100000111;
11'd363 : tab2 = 23'b01110001010001111001101;
11'd364 : tab2 = 23'b01110000111110010011111;
11'd365 : tab2 = 23'b01110000101010101111101;
11'd366 : tab2 = 23'b01110000010111001101001;
11'd367 : tab2 = 23'b01110000000011101100001;
11'd368 : tab2 = 23'b01101111110000001100101;
11'd369 : tab2 = 23'b01101111011100101110110;
11'd370 : tab2 = 23'b01101111001001010010011;
11'd371 : tab2 = 23'b01101110110101110111100;
11'd372 : tab2 = 23'b01101110100010011110011;
11'd373 : tab2 = 23'b01101110001111000110100;
11'd374 : tab2 = 23'b01101101111011110000011;
11'd375 : tab2 = 23'b01101101101000011011110;
11'd376 : tab2 = 23'b01101101010101001000100;
11'd377 : tab2 = 23'b01101101000001110110110;
11'd378 : tab2 = 23'b01101100101110100110110;
11'd379 : tab2 = 23'b01101100011011011000010;
11'd380 : tab2 = 23'b01101100001000001011001;
11'd381 : tab2 = 23'b01101011110100111111100;
11'd382 : tab2 = 23'b01101011100001110101011;
11'd383 : tab2 = 23'b01101011001110101100111;
11'd384 : tab2 = 23'b01101010111011100110000;
11'd385 : tab2 = 23'b01101010101000100000011;
11'd386 : tab2 = 23'b01101010010101011100100;
11'd387 : tab2 = 23'b01101010000010011010000;
11'd388 : tab2 = 23'b01101001101111011001001;
11'd389 : tab2 = 23'b01101001011100011001100;
11'd390 : tab2 = 23'b01101001001001011011101;
11'd391 : tab2 = 23'b01101000110110011111001;
11'd392 : tab2 = 23'b01101000100011100100000;
11'd393 : tab2 = 23'b01101000010000101010100;
11'd394 : tab2 = 23'b01100111111101110010100;
11'd395 : tab2 = 23'b01100111101010111011110;
11'd396 : tab2 = 23'b01100111011000000110101;
11'd397 : tab2 = 23'b01100111000101010011010;
11'd398 : tab2 = 23'b01100110110010100001001;
11'd399 : tab2 = 23'b01100110011111110000100;
11'd400 : tab2 = 23'b01100110001101000001010;
11'd401 : tab2 = 23'b01100101111010010011100;
11'd402 : tab2 = 23'b01100101100111100111010;
11'd403 : tab2 = 23'b01100101010100111100011;
11'd404 : tab2 = 23'b01100101000010010011001;
11'd405 : tab2 = 23'b01100100101111101011010;
11'd406 : tab2 = 23'b01100100011101000100110;
11'd407 : tab2 = 23'b01100100001010100000000;
11'd408 : tab2 = 23'b01100011110111111100011;
11'd409 : tab2 = 23'b01100011100101011010100;
11'd410 : tab2 = 23'b01100011010010111001101;
11'd411 : tab2 = 23'b01100011000000011010101;
11'd412 : tab2 = 23'b01100010101101111100110;
11'd413 : tab2 = 23'b01100010011011100000100;
11'd414 : tab2 = 23'b01100010001001000101101;
11'd415 : tab2 = 23'b01100001110110101100010;
11'd416 : tab2 = 23'b01100001100100010100011;
11'd417 : tab2 = 23'b01100001010001111101110;
11'd418 : tab2 = 23'b01100000111111101000101;
11'd419 : tab2 = 23'b01100000101101010101001;
11'd420 : tab2 = 23'b01100000011011000010111;
11'd421 : tab2 = 23'b01100000001000110001111;
11'd422 : tab2 = 23'b01011111110110100010100;
11'd423 : tab2 = 23'b01011111100100010100100;
11'd424 : tab2 = 23'b01011111010010000111111;
11'd425 : tab2 = 23'b01011110111111111100100;
11'd426 : tab2 = 23'b01011110101101110010111;
11'd427 : tab2 = 23'b01011110011011101010101;
11'd428 : tab2 = 23'b01011110001001100011110;
11'd429 : tab2 = 23'b01011101110111011110000;
11'd430 : tab2 = 23'b01011101100101011001110;
11'd431 : tab2 = 23'b01011101010011010111000;
11'd432 : tab2 = 23'b01011101000001010101111;
11'd433 : tab2 = 23'b01011100101111010101111;
11'd434 : tab2 = 23'b01011100011101010111010;
11'd435 : tab2 = 23'b01011100001011011010000;
11'd436 : tab2 = 23'b01011011111001011110001;
11'd437 : tab2 = 23'b01011011100111100011110;
11'd438 : tab2 = 23'b01011011010101101010111;
11'd439 : tab2 = 23'b01011011000011110011010;
11'd440 : tab2 = 23'b01011010110001111100110;
11'd441 : tab2 = 23'b01011010100000000111111;
11'd442 : tab2 = 23'b01011010001110010100011;
11'd443 : tab2 = 23'b01011001111100100010010;
11'd444 : tab2 = 23'b01011001101010110001100;
11'd445 : tab2 = 23'b01011001011001000010001;
11'd446 : tab2 = 23'b01011001000111010100001;
11'd447 : tab2 = 23'b01011000110101100111011;
11'd448 : tab2 = 23'b01011000100011111100001;
11'd449 : tab2 = 23'b01011000010010010010001;
11'd450 : tab2 = 23'b01011000000000101001100;
11'd451 : tab2 = 23'b01010111101111000010010;
11'd452 : tab2 = 23'b01010111011101011100010;
11'd453 : tab2 = 23'b01010111001011110111110;
11'd454 : tab2 = 23'b01010110111010010100100;
11'd455 : tab2 = 23'b01010110101000110010110;
11'd456 : tab2 = 23'b01010110010111010010010;
11'd457 : tab2 = 23'b01010110000101110011000;
11'd458 : tab2 = 23'b01010101110100010101010;
11'd459 : tab2 = 23'b01010101100010111000110;
11'd460 : tab2 = 23'b01010101010001011101101;
11'd461 : tab2 = 23'b01010101000000000011111;
11'd462 : tab2 = 23'b01010100101110101011011;
11'd463 : tab2 = 23'b01010100011101010100000;
11'd464 : tab2 = 23'b01010100001011111110010;
11'd465 : tab2 = 23'b01010011111010101001110;
11'd466 : tab2 = 23'b01010011101001010110101;
11'd467 : tab2 = 23'b01010011011000000100110;
11'd468 : tab2 = 23'b01010011000110110100001;
11'd469 : tab2 = 23'b01010010110101100100111;
11'd470 : tab2 = 23'b01010010100100010111000;
11'd471 : tab2 = 23'b01010010010011001010011;
11'd472 : tab2 = 23'b01010010000001111111001;
11'd473 : tab2 = 23'b01010001110000110100111;
11'd474 : tab2 = 23'b01010001011111101100011;
11'd475 : tab2 = 23'b01010001001110100100111;
11'd476 : tab2 = 23'b01010000111101011110111;
11'd477 : tab2 = 23'b01010000101100011010000;
11'd478 : tab2 = 23'b01010000011011010110110;
11'd479 : tab2 = 23'b01010000001010010100010;
11'd480 : tab2 = 23'b01001111111001010011011;
11'd481 : tab2 = 23'b01001111101000010011111;
11'd482 : tab2 = 23'b01001111010111010101100;
11'd483 : tab2 = 23'b01001111000110011000011;
11'd484 : tab2 = 23'b01001110110101011100110;
11'd485 : tab2 = 23'b01001110100100100010011;
11'd486 : tab2 = 23'b01001110010011101001000;
11'd487 : tab2 = 23'b01001110000010110001010;
11'd488 : tab2 = 23'b01001101110001111010110;
11'd489 : tab2 = 23'b01001101100001000101000;
11'd490 : tab2 = 23'b01001101010000010001000;
11'd491 : tab2 = 23'b01001100111111011110001;
11'd492 : tab2 = 23'b01001100101110101100110;
11'd493 : tab2 = 23'b01001100011101111100100;
11'd494 : tab2 = 23'b01001100001101001101100;
11'd495 : tab2 = 23'b01001011111100011111110;
11'd496 : tab2 = 23'b01001011101011110011011;
11'd497 : tab2 = 23'b01001011011011001000001;
11'd498 : tab2 = 23'b01001011001010011110000;
11'd499 : tab2 = 23'b01001010111001110101011;
11'd500 : tab2 = 23'b01001010101001001110000;
11'd501 : tab2 = 23'b01001010011000100111100;
11'd502 : tab2 = 23'b01001010001000000010100;
11'd503 : tab2 = 23'b01001001110111011111000;
11'd504 : tab2 = 23'b01001001100110111100100;
11'd505 : tab2 = 23'b01001001010110011011011;
11'd506 : tab2 = 23'b01001001000101111011011;
11'd507 : tab2 = 23'b01001000110101011100100;
11'd508 : tab2 = 23'b01001000100100111111000;
11'd509 : tab2 = 23'b01001000010100100010110;
11'd510 : tab2 = 23'b01001000000100000111110;
11'd511 : tab2 = 23'b01000111110011101110000;
11'd512 : tab2 = 23'b01000111100011010101011;
11'd513 : tab2 = 23'b01000111010010111110000;
11'd514 : tab2 = 23'b01000111000010101000000;
11'd515 : tab2 = 23'b01000110110010010011000;
11'd516 : tab2 = 23'b01000110100001111111010;
11'd517 : tab2 = 23'b01000110010001101100111;
11'd518 : tab2 = 23'b01000110000001011011110;
11'd519 : tab2 = 23'b01000101110001001011110;
11'd520 : tab2 = 23'b01000101100000111100101;
11'd521 : tab2 = 23'b01000101010000101111001;
11'd522 : tab2 = 23'b01000101000000100010110;
11'd523 : tab2 = 23'b01000100110000010111100;
11'd524 : tab2 = 23'b01000100100000001101101;
11'd525 : tab2 = 23'b01000100010000000100111;
11'd526 : tab2 = 23'b01000011111111111101010;
11'd527 : tab2 = 23'b01000011101111110110111;
11'd528 : tab2 = 23'b01000011011111110001110;
11'd529 : tab2 = 23'b01000011001111101101110;
11'd530 : tab2 = 23'b01000010111111101011000;
11'd531 : tab2 = 23'b01000010101111101001011;
11'd532 : tab2 = 23'b01000010011111101001000;
11'd533 : tab2 = 23'b01000010001111101001111;
11'd534 : tab2 = 23'b01000001111111101100000;
11'd535 : tab2 = 23'b01000001101111101111001;
11'd536 : tab2 = 23'b01000001011111110011100;
11'd537 : tab2 = 23'b01000001001111111001001;
11'd538 : tab2 = 23'b01000000111111111111110;
11'd539 : tab2 = 23'b01000000110000000111110;
11'd540 : tab2 = 23'b01000000100000010000111;
11'd541 : tab2 = 23'b01000000010000011011001;
11'd542 : tab2 = 23'b01000000000000100110011;
11'd543 : tab2 = 23'b00111111110000110011000;
11'd544 : tab2 = 23'b00111111100001000000111;
11'd545 : tab2 = 23'b00111111010001001111111;
11'd546 : tab2 = 23'b00111111000001100000000;
11'd547 : tab2 = 23'b00111110110001110001011;
11'd548 : tab2 = 23'b00111110100010000011110;
11'd549 : tab2 = 23'b00111110010010010111010;
11'd550 : tab2 = 23'b00111110000010101100001;
11'd551 : tab2 = 23'b00111101110011000010000;
11'd552 : tab2 = 23'b00111101100011011001000;
11'd553 : tab2 = 23'b00111101010011110001010;
11'd554 : tab2 = 23'b00111101000100001010101;
11'd555 : tab2 = 23'b00111100110100100101010;
11'd556 : tab2 = 23'b00111100100101000000111;
11'd557 : tab2 = 23'b00111100010101011101111;
11'd558 : tab2 = 23'b00111100000101111011101;
11'd559 : tab2 = 23'b00111011110110011010111;
11'd560 : tab2 = 23'b00111011100110111011001;
11'd561 : tab2 = 23'b00111011010111011100100;
11'd562 : tab2 = 23'b00111011000111111111000;
11'd563 : tab2 = 23'b00111010111000100010101;
11'd564 : tab2 = 23'b00111010101001000111100;
11'd565 : tab2 = 23'b00111010011001101101100;
11'd566 : tab2 = 23'b00111010001010010100110;
11'd567 : tab2 = 23'b00111001111010111100101;
11'd568 : tab2 = 23'b00111001101011100110001;
11'd569 : tab2 = 23'b00111001011100010000101;
11'd570 : tab2 = 23'b00111001001100111100010;
11'd571 : tab2 = 23'b00111000111101101000110;
11'd572 : tab2 = 23'b00111000101110010110110;
11'd573 : tab2 = 23'b00111000011111000101101;
11'd574 : tab2 = 23'b00111000001111110101111;
11'd575 : tab2 = 23'b00111000000000100111000;
11'd576 : tab2 = 23'b00110111110001011001000;
11'd577 : tab2 = 23'b00110111100010001100100;
11'd578 : tab2 = 23'b00110111010011000001001;
11'd579 : tab2 = 23'b00110111000011110110110;
11'd580 : tab2 = 23'b00110110110100101101100;
11'd581 : tab2 = 23'b00110110100101100101011;
11'd582 : tab2 = 23'b00110110010110011110010;
11'd583 : tab2 = 23'b00110110000111011000011;
11'd584 : tab2 = 23'b00110101111000010011100;
11'd585 : tab2 = 23'b00110101101001001111110;
11'd586 : tab2 = 23'b00110101011010001100111;
11'd587 : tab2 = 23'b00110101001011001011011;
11'd588 : tab2 = 23'b00110100111100001010111;
11'd589 : tab2 = 23'b00110100101101001011101;
11'd590 : tab2 = 23'b00110100011110001101001;
11'd591 : tab2 = 23'b00110100001111010000001;
11'd592 : tab2 = 23'b00110100000000010100000;
11'd593 : tab2 = 23'b00110011110001011000110;
11'd594 : tab2 = 23'b00110011100010011111000;
11'd595 : tab2 = 23'b00110011010011100110010;
11'd596 : tab2 = 23'b00110011000100101110010;
11'd597 : tab2 = 23'b00110010110101110111101;
11'd598 : tab2 = 23'b00110010100111000010001;
11'd599 : tab2 = 23'b00110010011000001101101;
11'd600 : tab2 = 23'b00110010001001011010001;
11'd601 : tab2 = 23'b00110001111010100111101;
11'd602 : tab2 = 23'b00110001101011110110010;
11'd603 : tab2 = 23'b00110001011101000110000;
11'd604 : tab2 = 23'b00110001001110010111000;
11'd605 : tab2 = 23'b00110000111111101000110;
11'd606 : tab2 = 23'b00110000110000111011110;
11'd607 : tab2 = 23'b00110000100010001111110;
11'd608 : tab2 = 23'b00110000010011100100101;
11'd609 : tab2 = 23'b00110000000100111011000;
11'd610 : tab2 = 23'b00101111110110010010000;
11'd611 : tab2 = 23'b00101111100111101010010;
11'd612 : tab2 = 23'b00101111011001000011100;
11'd613 : tab2 = 23'b00101111001010011110000;
11'd614 : tab2 = 23'b00101110111011111001010;
11'd615 : tab2 = 23'b00101110101101010101110;
11'd616 : tab2 = 23'b00101110011110110011010;
11'd617 : tab2 = 23'b00101110010000010001110;
11'd618 : tab2 = 23'b00101110000001110001011;
11'd619 : tab2 = 23'b00101101110011010010001;
11'd620 : tab2 = 23'b00101101100100110011110;
11'd621 : tab2 = 23'b00101101010110010110011;
11'd622 : tab2 = 23'b00101101000111111010010;
11'd623 : tab2 = 23'b00101100111001011111001;
11'd624 : tab2 = 23'b00101100101011000100111;
11'd625 : tab2 = 23'b00101100011100101011110;
11'd626 : tab2 = 23'b00101100001110010011100;
11'd627 : tab2 = 23'b00101011111111111100011;
11'd628 : tab2 = 23'b00101011110001100110011;
11'd629 : tab2 = 23'b00101011100011010001100;
11'd630 : tab2 = 23'b00101011010100111101100;
11'd631 : tab2 = 23'b00101011000110101010101;
11'd632 : tab2 = 23'b00101010111000011000110;
11'd633 : tab2 = 23'b00101010101010000111101;
11'd634 : tab2 = 23'b00101010011011110111110;
11'd635 : tab2 = 23'b00101010001101101000111;
11'd636 : tab2 = 23'b00101001111111011011001;
11'd637 : tab2 = 23'b00101001110001001110011;
11'd638 : tab2 = 23'b00101001100011000010011;
11'd639 : tab2 = 23'b00101001010100110111101;
11'd640 : tab2 = 23'b00101001000110101101101;
11'd641 : tab2 = 23'b00101000111000100100111;
11'd642 : tab2 = 23'b00101000101010011101001;
11'd643 : tab2 = 23'b00101000011100010110011;
11'd644 : tab2 = 23'b00101000001110010000101;
11'd645 : tab2 = 23'b00101000000000001011111;
11'd646 : tab2 = 23'b00100111110010001000001;
11'd647 : tab2 = 23'b00100111100100000101011;
11'd648 : tab2 = 23'b00100111010110000011101;
11'd649 : tab2 = 23'b00100111001000000010111;
11'd650 : tab2 = 23'b00100110111010000011001;
11'd651 : tab2 = 23'b00100110101100000100010;
11'd652 : tab2 = 23'b00100110011110000110101;
11'd653 : tab2 = 23'b00100110010000001001110;
11'd654 : tab2 = 23'b00100110000010001110000;
11'd655 : tab2 = 23'b00100101110100010011001;
11'd656 : tab2 = 23'b00100101100110011001011;
11'd657 : tab2 = 23'b00100101011000100000101;
11'd658 : tab2 = 23'b00100101001010101000110;
11'd659 : tab2 = 23'b00100100111100110001110;
11'd660 : tab2 = 23'b00100100101110111100000;
11'd661 : tab2 = 23'b00100100100001000111000;
11'd662 : tab2 = 23'b00100100010011010011000;
11'd663 : tab2 = 23'b00100100000101100000001;
11'd664 : tab2 = 23'b00100011110111101110010;
11'd665 : tab2 = 23'b00100011101001111101011;
11'd666 : tab2 = 23'b00100011011100001101010;
11'd667 : tab2 = 23'b00100011001110011110010;
11'd668 : tab2 = 23'b00100011000000110000010;
11'd669 : tab2 = 23'b00100010110011000011000;
11'd670 : tab2 = 23'b00100010100101010110111;
11'd671 : tab2 = 23'b00100010010111101011101;
11'd672 : tab2 = 23'b00100010001010000001100;
11'd673 : tab2 = 23'b00100001111100011000010;
11'd674 : tab2 = 23'b00100001101110110000000;
11'd675 : tab2 = 23'b00100001100001001000101;
11'd676 : tab2 = 23'b00100001010011100010010;
11'd677 : tab2 = 23'b00100001000101111100111;
11'd678 : tab2 = 23'b00100000111000011000011;
11'd679 : tab2 = 23'b00100000101010110101000;
11'd680 : tab2 = 23'b00100000011101010010011;
11'd681 : tab2 = 23'b00100000001111110001000;
11'd682 : tab2 = 23'b00100000000010010000010;
11'd683 : tab2 = 23'b00011111110100110000100;
11'd684 : tab2 = 23'b00011111100111010001101;
11'd685 : tab2 = 23'b00011111011001110011111;
11'd686 : tab2 = 23'b00011111001100010111010;
11'd687 : tab2 = 23'b00011110111110111011001;
11'd688 : tab2 = 23'b00011110110001100000010;
11'd689 : tab2 = 23'b00011110100100000110011;
11'd690 : tab2 = 23'b00011110010110101101001;
11'd691 : tab2 = 23'b00011110001001010101000;
11'd692 : tab2 = 23'b00011101111011111101111;
11'd693 : tab2 = 23'b00011101101110100111100;
11'd694 : tab2 = 23'b00011101100001010010010;
11'd695 : tab2 = 23'b00011101010011111101111;
11'd696 : tab2 = 23'b00011101000110101010011;
11'd697 : tab2 = 23'b00011100111001010111110;
11'd698 : tab2 = 23'b00011100101100000110011;
11'd699 : tab2 = 23'b00011100011110110101100;
11'd700 : tab2 = 23'b00011100010001100101110;
11'd701 : tab2 = 23'b00011100000100010110111;
11'd702 : tab2 = 23'b00011011110111001001001;
11'd703 : tab2 = 23'b00011011101001111100001;
11'd704 : tab2 = 23'b00011011011100110000000;
11'd705 : tab2 = 23'b00011011001111100101000;
11'd706 : tab2 = 23'b00011011000010011010101;
11'd707 : tab2 = 23'b00011010110101010001010;
11'd708 : tab2 = 23'b00011010101000001000111;
11'd709 : tab2 = 23'b00011010011011000001100;
11'd710 : tab2 = 23'b00011010001101111010111;
11'd711 : tab2 = 23'b00011010000000110101011;
11'd712 : tab2 = 23'b00011001110011110000101;
11'd713 : tab2 = 23'b00011001100110101100110;
11'd714 : tab2 = 23'b00011001011001101001111;
11'd715 : tab2 = 23'b00011001001100100111101;
11'd716 : tab2 = 23'b00011000111111100110101;
11'd717 : tab2 = 23'b00011000110010100110010;
11'd718 : tab2 = 23'b00011000100101100111001;
11'd719 : tab2 = 23'b00011000011000101000110;
11'd720 : tab2 = 23'b00011000001011101011001;
11'd721 : tab2 = 23'b00010111111110101110100;
11'd722 : tab2 = 23'b00010111110001110010111;
11'd723 : tab2 = 23'b00010111100100111000000;
11'd724 : tab2 = 23'b00010111010111111110010;
11'd725 : tab2 = 23'b00010111001011000101000;
11'd726 : tab2 = 23'b00010110111110001100111;
11'd727 : tab2 = 23'b00010110110001010101101;
11'd728 : tab2 = 23'b00010110100100011111010;
11'd729 : tab2 = 23'b00010110010111101001111;
11'd730 : tab2 = 23'b00010110001010110101011;
11'd731 : tab2 = 23'b00010101111110000001100;
11'd732 : tab2 = 23'b00010101110001001110101;
11'd733 : tab2 = 23'b00010101100100011100111;
11'd734 : tab2 = 23'b00010101010111101011110;
11'd735 : tab2 = 23'b00010101001010111011101;
11'd736 : tab2 = 23'b00010100111110001100011;
11'd737 : tab2 = 23'b00010100110001011101110;
11'd738 : tab2 = 23'b00010100100100110000011;
11'd739 : tab2 = 23'b00010100011000000011101;
11'd740 : tab2 = 23'b00010100001011010111111;
11'd741 : tab2 = 23'b00010011111110101100111;
11'd742 : tab2 = 23'b00010011110010000010111;
11'd743 : tab2 = 23'b00010011100101011001111;
11'd744 : tab2 = 23'b00010011011000110001100;
11'd745 : tab2 = 23'b00010011001100001010000;
11'd746 : tab2 = 23'b00010010111111100011100;
11'd747 : tab2 = 23'b00010010110010111101111;
11'd748 : tab2 = 23'b00010010100110011000111;
11'd749 : tab2 = 23'b00010010011001110100111;
11'd750 : tab2 = 23'b00010010001101010010000;
11'd751 : tab2 = 23'b00010010000000101111101;
11'd752 : tab2 = 23'b00010001110100001110010;
11'd753 : tab2 = 23'b00010001100111101101110;
11'd754 : tab2 = 23'b00010001011011001110000;
11'd755 : tab2 = 23'b00010001001110101111001;
11'd756 : tab2 = 23'b00010001000010010001010;
11'd757 : tab2 = 23'b00010000110101110100001;
11'd758 : tab2 = 23'b00010000101001010111111;
11'd759 : tab2 = 23'b00010000011100111100011;
11'd760 : tab2 = 23'b00010000010000100001110;
11'd761 : tab2 = 23'b00010000000100001000001;
11'd762 : tab2 = 23'b00001111110111101111010;
11'd763 : tab2 = 23'b00001111101011010111010;
11'd764 : tab2 = 23'b00001111011110111111111;
11'd765 : tab2 = 23'b00001111010010101001101;
11'd766 : tab2 = 23'b00001111000110010100011;
11'd767 : tab2 = 23'b00001110111001111111110;
11'd768 : tab2 = 23'b00001110101101101011110;
11'd769 : tab2 = 23'b00001110100001011000110;
11'd770 : tab2 = 23'b00001110010101000110110;
11'd771 : tab2 = 23'b00001110001000110101011;
11'd772 : tab2 = 23'b00001101111100100100111;
11'd773 : tab2 = 23'b00001101110000010101011;
11'd774 : tab2 = 23'b00001101100100000110100;
11'd775 : tab2 = 23'b00001101010111111000101;
11'd776 : tab2 = 23'b00001101001011101011011;
11'd777 : tab2 = 23'b00001100111111011111001;
11'd778 : tab2 = 23'b00001100110011010011110;
11'd779 : tab2 = 23'b00001100100111001000111;
11'd780 : tab2 = 23'b00001100011010111111001;
11'd781 : tab2 = 23'b00001100001110110110000;
11'd782 : tab2 = 23'b00001100000010101101111;
11'd783 : tab2 = 23'b00001011110110100110110;
11'd784 : tab2 = 23'b00001011101010100000000;
11'd785 : tab2 = 23'b00001011011110011010011;
11'd786 : tab2 = 23'b00001011010010010101100;
11'd787 : tab2 = 23'b00001011000110010001011;
11'd788 : tab2 = 23'b00001010111010001110001;
11'd789 : tab2 = 23'b00001010101110001011110;
11'd790 : tab2 = 23'b00001010100010001010001;
11'd791 : tab2 = 23'b00001010010110001001001;
11'd792 : tab2 = 23'b00001010001010001001001;
11'd793 : tab2 = 23'b00001001111110001010001;
11'd794 : tab2 = 23'b00001001110010001011110;
11'd795 : tab2 = 23'b00001001100110001110000;
11'd796 : tab2 = 23'b00001001011010010001010;
11'd797 : tab2 = 23'b00001001001110010101011;
11'd798 : tab2 = 23'b00001001000010011010010;
11'd799 : tab2 = 23'b00001000110110011111110;
11'd800 : tab2 = 23'b00001000101010100110010;
11'd801 : tab2 = 23'b00001000011110101101100;
11'd802 : tab2 = 23'b00001000010010110101101;
11'd803 : tab2 = 23'b00001000000110111110100;
11'd804 : tab2 = 23'b00000111111011001000000;
11'd805 : tab2 = 23'b00000111101111010010100;
11'd806 : tab2 = 23'b00000111100011011101111;
11'd807 : tab2 = 23'b00000111010111101001110;
11'd808 : tab2 = 23'b00000111001011110110101;
11'd809 : tab2 = 23'b00000111000000000100001;
11'd810 : tab2 = 23'b00000110110100010010110;
11'd811 : tab2 = 23'b00000110101000100001111;
11'd812 : tab2 = 23'b00000110011100110001111;
11'd813 : tab2 = 23'b00000110010001000010101;
11'd814 : tab2 = 23'b00000110000101010100010;
11'd815 : tab2 = 23'b00000101111001100110100;
11'd816 : tab2 = 23'b00000101101101111001101;
11'd817 : tab2 = 23'b00000101100010001101101;
11'd818 : tab2 = 23'b00000101010110100010010;
11'd819 : tab2 = 23'b00000101001010110111111;
11'd820 : tab2 = 23'b00000100111111001110001;
11'd821 : tab2 = 23'b00000100110011100101001;
11'd822 : tab2 = 23'b00000100100111111101000;
11'd823 : tab2 = 23'b00000100011100010101100;
11'd824 : tab2 = 23'b00000100010000101111000;
11'd825 : tab2 = 23'b00000100000101001001001;
11'd826 : tab2 = 23'b00000011111001100100000;
11'd827 : tab2 = 23'b00000011101101111111110;
11'd828 : tab2 = 23'b00000011100010011100001;
11'd829 : tab2 = 23'b00000011010110111001100;
11'd830 : tab2 = 23'b00000011001011010111100;
11'd831 : tab2 = 23'b00000010111111110110011;
11'd832 : tab2 = 23'b00000010110100010101111;
11'd833 : tab2 = 23'b00000010101000110110001;
11'd834 : tab2 = 23'b00000010011101010111001;
11'd835 : tab2 = 23'b00000010010001111001000;
11'd836 : tab2 = 23'b00000010000110011011110;
11'd837 : tab2 = 23'b00000001111010111111000;
11'd838 : tab2 = 23'b00000001101111100011001;
11'd839 : tab2 = 23'b00000001100100001000000;
11'd840 : tab2 = 23'b00000001011000101101110;
11'd841 : tab2 = 23'b00000001001101010100001;
11'd842 : tab2 = 23'b00000001000001111011010;
11'd843 : tab2 = 23'b00000000110110100011010;
11'd844 : tab2 = 23'b00000000101011001011111;
11'd845 : tab2 = 23'b00000000011111110101010;
11'd846 : tab2 = 23'b00000000010100011111100;
11'd847 : tab2 = 23'b00000000001001001010011;
11'd848 : tab2 = 23'b11111111111011101100100;
11'd849 : tab2 = 23'b11111111100101000101001;
11'd850 : tab2 = 23'b11111111001110011111100;
11'd851 : tab2 = 23'b11111110110111111011100;
11'd852 : tab2 = 23'b11111110100001011000110;
11'd853 : tab2 = 23'b11111110001010110111100;
11'd854 : tab2 = 23'b11111101110100011000010;
11'd855 : tab2 = 23'b11111101011101111001110;
11'd856 : tab2 = 23'b11111101000111011101001;
11'd857 : tab2 = 23'b11111100110001000001111;
11'd858 : tab2 = 23'b11111100011010101000011;
11'd859 : tab2 = 23'b11111100000100010000001;
11'd860 : tab2 = 23'b11111011101101111001000;
11'd861 : tab2 = 23'b11111011010111100011111;
11'd862 : tab2 = 23'b11111011000001001111111;
11'd863 : tab2 = 23'b11111010101010111101111;
11'd864 : tab2 = 23'b11111010010100101101000;
11'd865 : tab2 = 23'b11111001111110011101010;
11'd866 : tab2 = 23'b11111001101000001111100;
11'd867 : tab2 = 23'b11111001010010000010111;
11'd868 : tab2 = 23'b11111000111011111000001;
11'd869 : tab2 = 23'b11111000100101101110101;
11'd870 : tab2 = 23'b11111000001111100110010;
11'd871 : tab2 = 23'b11110111111001011111111;
11'd872 : tab2 = 23'b11110111100011011010101;
11'd873 : tab2 = 23'b11110111001101010110111;
11'd874 : tab2 = 23'b11110110110111010100101;
11'd875 : tab2 = 23'b11110110100001010011101;
11'd876 : tab2 = 23'b11110110001011010100010;
11'd877 : tab2 = 23'b11110101110101010110010;
11'd878 : tab2 = 23'b11110101011111011001100;
11'd879 : tab2 = 23'b11110101001001011110101;
11'd880 : tab2 = 23'b11110100110011100100111;
11'd881 : tab2 = 23'b11110100011101101101001;
11'd882 : tab2 = 23'b11110100000111110110001;
11'd883 : tab2 = 23'b11110011110010000001000;
11'd884 : tab2 = 23'b11110011011100001100101;
11'd885 : tab2 = 23'b11110011000110011010010;
11'd886 : tab2 = 23'b11110010110000101001010;
11'd887 : tab2 = 23'b11110010011010111001101;
11'd888 : tab2 = 23'b11110010000101001011011;
11'd889 : tab2 = 23'b11110001101111011111000;
11'd890 : tab2 = 23'b11110001011001110011001;
11'd891 : tab2 = 23'b11110001000100001001001;
11'd892 : tab2 = 23'b11110000101110100001000;
11'd893 : tab2 = 23'b11110000011000111001101;
11'd894 : tab2 = 23'b11110000000011010011111;
11'd895 : tab2 = 23'b11101111101101101111101;
11'd896 : tab2 = 23'b11101111011000001100110;
11'd897 : tab2 = 23'b11101111000010101011001;
11'd898 : tab2 = 23'b11101110101101001011001;
11'd899 : tab2 = 23'b11101110010111101100100;
11'd900 : tab2 = 23'b11101110000010001111011;
11'd901 : tab2 = 23'b11101101101100110011001;
11'd902 : tab2 = 23'b11101101010111011000101;
11'd903 : tab2 = 23'b11101101000001111111011;
11'd904 : tab2 = 23'b11101100101100101000000;
11'd905 : tab2 = 23'b11101100010111010001011;
11'd906 : tab2 = 23'b11101100000001111100101;
11'd907 : tab2 = 23'b11101011101100101000101;
11'd908 : tab2 = 23'b11101011010111010110101;
11'd909 : tab2 = 23'b11101011000010000110000;
11'd910 : tab2 = 23'b11101010101100110110100;
11'd911 : tab2 = 23'b11101010010111101000101;
11'd912 : tab2 = 23'b11101010000010011011110;
11'd913 : tab2 = 23'b11101001101101010000100;
11'd914 : tab2 = 23'b11101001011000000110101;
11'd915 : tab2 = 23'b11101001000010111110000;
11'd916 : tab2 = 23'b11101000101101110110111;
11'd917 : tab2 = 23'b11101000011000110001001;
11'd918 : tab2 = 23'b11101000000011101100101;
11'd919 : tab2 = 23'b11100111101110101001010;
11'd920 : tab2 = 23'b11100111011001100111110;
11'd921 : tab2 = 23'b11100111000100100111010;
11'd922 : tab2 = 23'b11100110101111101000000;
11'd923 : tab2 = 23'b11100110011010101010101;
11'd924 : tab2 = 23'b11100110000101101110010;
11'd925 : tab2 = 23'b11100101110000110011001;
11'd926 : tab2 = 23'b11100101011011111001110;
11'd927 : tab2 = 23'b11100101000111000001101;
11'd928 : tab2 = 23'b11100100110010001010100;
11'd929 : tab2 = 23'b11100100011101010101011;
11'd930 : tab2 = 23'b11100100001000100000111;
11'd931 : tab2 = 23'b11100011110011101101111;
11'd932 : tab2 = 23'b11100011011110111100100;
11'd933 : tab2 = 23'b11100011001010001100011;
11'd934 : tab2 = 23'b11100010110101011101100;
11'd935 : tab2 = 23'b11100010100000101111111;
11'd936 : tab2 = 23'b11100010001100000011111;
11'd937 : tab2 = 23'b11100001110111011000110;
11'd938 : tab2 = 23'b11100001100010101111011;
11'd939 : tab2 = 23'b11100001001110000110111;
11'd940 : tab2 = 23'b11100000111001100000001;
11'd941 : tab2 = 23'b11100000100100111010101;
11'd942 : tab2 = 23'b11100000010000010110001;
11'd943 : tab2 = 23'b11011111111011110011011;
11'd944 : tab2 = 23'b11011111100111010001111;
11'd945 : tab2 = 23'b11011111010010110001100;
11'd946 : tab2 = 23'b11011110111110010010111;
11'd947 : tab2 = 23'b11011110101001110100110;
11'd948 : tab2 = 23'b11011110010101011000101;
11'd949 : tab2 = 23'b11011110000000111101110;
11'd950 : tab2 = 23'b11011101101100100011101;
11'd951 : tab2 = 23'b11011101011000001011010;
11'd952 : tab2 = 23'b11011101000011110100001;
11'd953 : tab2 = 23'b11011100101111011110101;
11'd954 : tab2 = 23'b11011100011011001001110;
11'd955 : tab2 = 23'b11011100000110110110100;
11'd956 : tab2 = 23'b11011011110010100100100;
11'd957 : tab2 = 23'b11011011011110010100001;
11'd958 : tab2 = 23'b11011011001010000100101;
11'd959 : tab2 = 23'b11011010110101110110101;
11'd960 : tab2 = 23'b11011010100001101010000;
11'd961 : tab2 = 23'b11011010001101011110010;
11'd962 : tab2 = 23'b11011001111001010100001;
11'd963 : tab2 = 23'b11011001100101001011010;
11'd964 : tab2 = 23'b11011001010001000011110;
11'd965 : tab2 = 23'b11011000111100111101011;
11'd966 : tab2 = 23'b11011000101000111000100;
11'd967 : tab2 = 23'b11011000010100110100101;
11'd968 : tab2 = 23'b11011000000000110001111;
11'd969 : tab2 = 23'b11010111101100110001000;
11'd970 : tab2 = 23'b11010111011000110001001;
11'd971 : tab2 = 23'b11010111000100110010011;
11'd972 : tab2 = 23'b11010110110000110100110;
11'd973 : tab2 = 23'b11010110011100111001000;
11'd974 : tab2 = 23'b11010110001000111101111;
11'd975 : tab2 = 23'b11010101110101000100010;
11'd976 : tab2 = 23'b11010101100001001100000;
11'd977 : tab2 = 23'b11010101001101010100101;
11'd978 : tab2 = 23'b11010100111001011110111;
11'd979 : tab2 = 23'b11010100100101101010010;
11'd980 : tab2 = 23'b11010100010001110111001;
11'd981 : tab2 = 23'b11010011111110000101001;
11'd982 : tab2 = 23'b11010011101010010100100;
11'd983 : tab2 = 23'b11010011010110100100101;
11'd984 : tab2 = 23'b11010011000010110110100;
11'd985 : tab2 = 23'b11010010101111001001001;
11'd986 : tab2 = 23'b11010010011011011101101;
11'd987 : tab2 = 23'b11010010000111110011001;
11'd988 : tab2 = 23'b11010001110100001001101;
11'd989 : tab2 = 23'b11010001100000100001011;
11'd990 : tab2 = 23'b11010001001100111010111;
11'd991 : tab2 = 23'b11010000111001010101011;
11'd992 : tab2 = 23'b11010000100101110001000;
11'd993 : tab2 = 23'b11010000010010001101101;
11'd994 : tab2 = 23'b11001111111110101100001;
11'd995 : tab2 = 23'b11001111101011001011000;
11'd996 : tab2 = 23'b11001111010111101011101;
11'd997 : tab2 = 23'b11001111000100001101011;
11'd998 : tab2 = 23'b11001110110000110000111;
11'd999 : tab2 = 23'b11001110011101010100110;
11'd1000 : tab2 = 23'b11001110001001111010011;
11'd1001 : tab2 = 23'b11001101110110100001000;
11'd1002 : tab2 = 23'b11001101100011001000111;
11'd1003 : tab2 = 23'b11001101001111110010011;
11'd1004 : tab2 = 23'b11001100111100011100010;
11'd1005 : tab2 = 23'b11001100101001001000000;
11'd1006 : tab2 = 23'b11001100010101110100110;
11'd1007 : tab2 = 23'b11001100000010100010101;
11'd1008 : tab2 = 23'b11001011101111010010001;
11'd1009 : tab2 = 23'b11001011011100000010001;
11'd1010 : tab2 = 23'b11001011001000110011111;
11'd1011 : tab2 = 23'b11001010110101100110101;
11'd1012 : tab2 = 23'b11001010100010011010111;
11'd1013 : tab2 = 23'b11001010001111010000001;
11'd1014 : tab2 = 23'b11001001111100000110100;
11'd1015 : tab2 = 23'b11001001101000111110010;
11'd1016 : tab2 = 23'b11001001010101110111000;
11'd1017 : tab2 = 23'b11001001000010110001010;
11'd1018 : tab2 = 23'b11001000101111101100010;
11'd1019 : tab2 = 23'b11001000011100101000111;
11'd1020 : tab2 = 23'b11001000001001100110011;
11'd1021 : tab2 = 23'b11000111110110100101001;
11'd1022 : tab2 = 23'b11000111100011100101011;
11'd1023 : tab2 = 23'b11000111010000100110010;
11'd1024 : tab2 = 23'b11000110111101101001000;
11'd1025 : tab2 = 23'b11000110101010101100011;
11'd1026 : tab2 = 23'b11000110010111110001001;
11'd1027 : tab2 = 23'b11000110000100110111000;
11'd1028 : tab2 = 23'b11000101110001111110010;
11'd1029 : tab2 = 23'b11000101011111000110001;
11'd1030 : tab2 = 23'b11000101001100001111111;
11'd1031 : tab2 = 23'b11000100111001011010010;
11'd1032 : tab2 = 23'b11000100100110100110001;
11'd1033 : tab2 = 23'b11000100010011110011010;
11'd1034 : tab2 = 23'b11000100000001000001001;
11'd1035 : tab2 = 23'b11000011101110010000111;
11'd1036 : tab2 = 23'b11000011011011100000111;
11'd1037 : tab2 = 23'b11000011001000110010101;
11'd1038 : tab2 = 23'b11000010110110000101011;
11'd1039 : tab2 = 23'b11000010100011011001100;
11'd1040 : tab2 = 23'b11000010010000101110110;
11'd1041 : tab2 = 23'b11000001111110000100110;
11'd1042 : tab2 = 23'b11000001101011011100011;
11'd1043 : tab2 = 23'b11000001011000110101000;
11'd1044 : tab2 = 23'b11000001000110001110110;
11'd1045 : tab2 = 23'b11000000110011101001101;
11'd1046 : tab2 = 23'b11000000100001000101110;
11'd1047 : tab2 = 23'b11000000001110100011000;
11'd1048 : tab2 = 23'b10111111111100000001101;
11'd1049 : tab2 = 23'b10111111101001100000111;
11'd1050 : tab2 = 23'b10111111010111000001101;
11'd1051 : tab2 = 23'b10111111000100100011010;
11'd1052 : tab2 = 23'b10111110110010000110011;
11'd1053 : tab2 = 23'b10111110011111101010010;
11'd1054 : tab2 = 23'b10111110001101001111110;
11'd1055 : tab2 = 23'b10111101111010110110010;
11'd1056 : tab2 = 23'b10111101101000011101100;
11'd1057 : tab2 = 23'b10111101010110000110001;
11'd1058 : tab2 = 23'b10111101000011110000001;
11'd1059 : tab2 = 23'b10111100110001011010111;
11'd1060 : tab2 = 23'b10111100011111000111010;
11'd1061 : tab2 = 23'b10111100001100110100000;
11'd1062 : tab2 = 23'b10111011111010100010100;
11'd1063 : tab2 = 23'b10111011101000010010000;
11'd1064 : tab2 = 23'b10111011010110000010100;
11'd1065 : tab2 = 23'b10111011000011110100001;
11'd1066 : tab2 = 23'b10111010110001100111000;
11'd1067 : tab2 = 23'b10111010011111011011000;
11'd1068 : tab2 = 23'b10111010001101010000010;
11'd1069 : tab2 = 23'b10111001111011000110000;
11'd1070 : tab2 = 23'b10111001101000111101011;
11'd1071 : tab2 = 23'b10111001010110110110001;
11'd1072 : tab2 = 23'b10111001000100101111100;
11'd1073 : tab2 = 23'b10111000110010101010011;
11'd1074 : tab2 = 23'b10111000100000100101110;
11'd1075 : tab2 = 23'b10111000001110100011000;
11'd1076 : tab2 = 23'b10110111111100100000100;
11'd1077 : tab2 = 23'b10110111101010011111110;
11'd1078 : tab2 = 23'b10110111011000100000000;
11'd1079 : tab2 = 23'b10110111000110100001010;
11'd1080 : tab2 = 23'b10110110110100100011100;
11'd1081 : tab2 = 23'b10110110100010100111010;
11'd1082 : tab2 = 23'b10110110010000101011111;
11'd1083 : tab2 = 23'b10110101111110110001010;
11'd1084 : tab2 = 23'b10110101101100111000010;
11'd1085 : tab2 = 23'b10110101011011000000010;
11'd1086 : tab2 = 23'b10110101001001001001000;
11'd1087 : tab2 = 23'b10110100110111010011001;
11'd1088 : tab2 = 23'b10110100100101011110010;
11'd1089 : tab2 = 23'b10110100010011101010101;
11'd1090 : tab2 = 23'b10110100000001110111110;
11'd1091 : tab2 = 23'b10110011110000000110101;
11'd1092 : tab2 = 23'b10110011011110010101110;
11'd1093 : tab2 = 23'b10110011001100100110101;
11'd1094 : tab2 = 23'b10110010111010111000001;
11'd1095 : tab2 = 23'b10110010101001001011000;
11'd1096 : tab2 = 23'b10110010010111011110111;
11'd1097 : tab2 = 23'b10110010000101110011110;
11'd1098 : tab2 = 23'b10110001110100001001111;
11'd1099 : tab2 = 23'b10110001100010100000111;
11'd1100 : tab2 = 23'b10110001010000111000110;
11'd1101 : tab2 = 23'b10110000111111010010010;
11'd1102 : tab2 = 23'b10110000101101101100100;
11'd1103 : tab2 = 23'b10110000011100000111110;
11'd1104 : tab2 = 23'b10110000001010100100011;
11'd1105 : tab2 = 23'b10101111111001000010000;
11'd1106 : tab2 = 23'b10101111100111100000101;
11'd1107 : tab2 = 23'b10101111010110000000010;
11'd1108 : tab2 = 23'b10101111000100100000110;
11'd1109 : tab2 = 23'b10101110110011000010110;
11'd1110 : tab2 = 23'b10101110100001100101101;
11'd1111 : tab2 = 23'b10101110010000001001010;
11'd1112 : tab2 = 23'b10101101111110101110100;
11'd1113 : tab2 = 23'b10101101101101010100001;
11'd1114 : tab2 = 23'b10101101011011111011100;
11'd1115 : tab2 = 23'b10101101001010100011110;
11'd1116 : tab2 = 23'b10101100111001001101000;
11'd1117 : tab2 = 23'b10101100100111110110111;
11'd1118 : tab2 = 23'b10101100010110100010001;
11'd1119 : tab2 = 23'b10101100000101001110110;
11'd1120 : tab2 = 23'b10101011110011111100000;
11'd1121 : tab2 = 23'b10101011100010101010101;
11'd1122 : tab2 = 23'b10101011010001011010001;
11'd1123 : tab2 = 23'b10101011000000001010011;
11'd1124 : tab2 = 23'b10101010101110111100010;
11'd1125 : tab2 = 23'b10101010011101101110100;
11'd1126 : tab2 = 23'b10101010001100100010011;
11'd1127 : tab2 = 23'b10101001111011010111010;
11'd1128 : tab2 = 23'b10101001101010001100110;
11'd1129 : tab2 = 23'b10101001011001000011100;
11'd1130 : tab2 = 23'b10101001000111111011011;
11'd1131 : tab2 = 23'b10101000110110110100001;
11'd1132 : tab2 = 23'b10101000100101101110000;
11'd1133 : tab2 = 23'b10101000010100101001001;
11'd1134 : tab2 = 23'b10101000000011100100111;
11'd1135 : tab2 = 23'b10100111110010100001101;
11'd1136 : tab2 = 23'b10100111100001100000000;
11'd1137 : tab2 = 23'b10100111010000011110110;
11'd1138 : tab2 = 23'b10100110111111011111001;
11'd1139 : tab2 = 23'b10100110101110011111111;
11'd1140 : tab2 = 23'b10100110011101100010001;
11'd1141 : tab2 = 23'b10100110001100100101001;
11'd1142 : tab2 = 23'b10100101111011101001001;
11'd1143 : tab2 = 23'b10100101101010101110011;
11'd1144 : tab2 = 23'b10100101011001110100101;
11'd1145 : tab2 = 23'b10100101001000111011111;
11'd1146 : tab2 = 23'b10100100111000000100001;
11'd1147 : tab2 = 23'b10100100100111001101010;
11'd1148 : tab2 = 23'b10100100010110010111100;
11'd1149 : tab2 = 23'b10100100000101100010101;
11'd1150 : tab2 = 23'b10100011110100101110110;
11'd1151 : tab2 = 23'b10100011100011111100001;
11'd1152 : tab2 = 23'b10100011010011001010101;
11'd1153 : tab2 = 23'b10100011000010011001101;
11'd1154 : tab2 = 23'b10100010110001101010000;
11'd1155 : tab2 = 23'b10100010100000111011010;
11'd1156 : tab2 = 23'b10100010010000001101010;
11'd1157 : tab2 = 23'b10100001111111100000111;
11'd1158 : tab2 = 23'b10100001101110110100110;
11'd1159 : tab2 = 23'b10100001011110001010011;
11'd1160 : tab2 = 23'b10100001001101100000111;
11'd1161 : tab2 = 23'b10100000111100110111101;
11'd1162 : tab2 = 23'b10100000101100010000001;
11'd1163 : tab2 = 23'b10100000011011101001100;
11'd1164 : tab2 = 23'b10100000001011000011101;
11'd1165 : tab2 = 23'b10011111111010011110101;
11'd1166 : tab2 = 23'b10011111101001111010111;
11'd1167 : tab2 = 23'b10011111011001011000010;
11'd1168 : tab2 = 23'b10011111001000110110100;
11'd1169 : tab2 = 23'b10011110111000010101101;
11'd1170 : tab2 = 23'b10011110100111110101111;
11'd1171 : tab2 = 23'b10011110010111010111000;
11'd1172 : tab2 = 23'b10011110000110111001001;
11'd1173 : tab2 = 23'b10011101110110011100001;
11'd1174 : tab2 = 23'b10011101100110000000100;
11'd1175 : tab2 = 23'b10011101010101100101100;
11'd1176 : tab2 = 23'b10011101000101001011100;
11'd1177 : tab2 = 23'b10011100110100110010110;
11'd1178 : tab2 = 23'b10011100100100011010101;
11'd1179 : tab2 = 23'b10011100010100000011011;
11'd1180 : tab2 = 23'b10011100000011101101100;
11'd1181 : tab2 = 23'b10011011110011011000101;
11'd1182 : tab2 = 23'b10011011100011000100010;
11'd1183 : tab2 = 23'b10011011010010110001010;
11'd1184 : tab2 = 23'b10011011000010011111010;
11'd1185 : tab2 = 23'b10011010110010001101110;
11'd1186 : tab2 = 23'b10011010100001111101101;
11'd1187 : tab2 = 23'b10011010010001101110100;
11'd1188 : tab2 = 23'b10011010000001011111111;
11'd1189 : tab2 = 23'b10011001110001010010111;
11'd1190 : tab2 = 23'b10011001100001000110010;
11'd1191 : tab2 = 23'b10011001010000111010111;
11'd1192 : tab2 = 23'b10011001000000110000100;
11'd1193 : tab2 = 23'b10011000110000100110101;
11'd1194 : tab2 = 23'b10011000100000011110100;
11'd1195 : tab2 = 23'b10011000010000010110101;
11'd1196 : tab2 = 23'b10011000000000010000010;
11'd1197 : tab2 = 23'b10010111110000001010010;
11'd1198 : tab2 = 23'b10010111100000000101111;
11'd1199 : tab2 = 23'b10010111010000000001110;
11'd1200 : tab2 = 23'b10010110111111111111010;
11'd1201 : tab2 = 23'b10010110101111111101000;
11'd1202 : tab2 = 23'b10010110011111111100011;
11'd1203 : tab2 = 23'b10010110001111111100001;
11'd1204 : tab2 = 23'b10010101111111111101011;
11'd1205 : tab2 = 23'b10010101101111111110111;
11'd1206 : tab2 = 23'b10010101100000000010000;
11'd1207 : tab2 = 23'b10010101010000000101100;
11'd1208 : tab2 = 23'b10010101000000001010100;
11'd1209 : tab2 = 23'b10010100110000001111111;
11'd1210 : tab2 = 23'b10010100100000010110110;
11'd1211 : tab2 = 23'b10010100010000011110000;
11'd1212 : tab2 = 23'b10010100000000100110111;
11'd1213 : tab2 = 23'b10010011110000101111111;
11'd1214 : tab2 = 23'b10010011100000111010101;
11'd1215 : tab2 = 23'b10010011010001000101101;
11'd1216 : tab2 = 23'b10010011000001010001111;
11'd1217 : tab2 = 23'b10010010110001011111000;
11'd1218 : tab2 = 23'b10010010100001101100110;
11'd1219 : tab2 = 23'b10010010010001111100001;
11'd1220 : tab2 = 23'b10010010000010001011111;
11'd1221 : tab2 = 23'b10010001110010011100110;
11'd1222 : tab2 = 23'b10010001100010101110101;
11'd1223 : tab2 = 23'b10010001010011000001000;
11'd1224 : tab2 = 23'b10010001000011010100110;
11'd1225 : tab2 = 23'b10010000110011101001001;
11'd1226 : tab2 = 23'b10010000100011111110101;
11'd1227 : tab2 = 23'b10010000010100010100111;
11'd1228 : tab2 = 23'b10010000000100101100011;
11'd1229 : tab2 = 23'b10001111110101000100011;
11'd1230 : tab2 = 23'b10001111100101011101110;
11'd1231 : tab2 = 23'b10001111010101110111101;
11'd1232 : tab2 = 23'b10001111000110010010100;
11'd1233 : tab2 = 23'b10001110110110101110010;
11'd1234 : tab2 = 23'b10001110100111001011000;
11'd1235 : tab2 = 23'b10001110010111101000101;
11'd1236 : tab2 = 23'b10001110001000000111001;
11'd1237 : tab2 = 23'b10001101111000100110101;
11'd1238 : tab2 = 23'b10001101101001000111000;
11'd1239 : tab2 = 23'b10001101011001101000011;
11'd1240 : tab2 = 23'b10001101001010001010101;
11'd1241 : tab2 = 23'b10001100111010101101110;
11'd1242 : tab2 = 23'b10001100101011010001101;
11'd1243 : tab2 = 23'b10001100011011110110010;
11'd1244 : tab2 = 23'b10001100001100011100010;
11'd1245 : tab2 = 23'b10001011111101000011001;
11'd1246 : tab2 = 23'b10001011101101101010010;
11'd1247 : tab2 = 23'b10001011011110010011000;
11'd1248 : tab2 = 23'b10001011001110111100101;
11'd1249 : tab2 = 23'b10001010111111100110101;
11'd1250 : tab2 = 23'b10001010110000010010000;
11'd1251 : tab2 = 23'b10001010100000111101110;
11'd1252 : tab2 = 23'b10001010010001101010110;
11'd1253 : tab2 = 23'b10001010000010011000110;
11'd1254 : tab2 = 23'b10001001110011000111010;
11'd1255 : tab2 = 23'b10001001100011110111000;
11'd1256 : tab2 = 23'b10001001010100100111101;
11'd1257 : tab2 = 23'b10001001000101011000111;
11'd1258 : tab2 = 23'b10001000110110001011001;
11'd1259 : tab2 = 23'b10001000100110111110001;
11'd1260 : tab2 = 23'b10001000010111110010001;
11'd1261 : tab2 = 23'b10001000001000100111001;
11'd1262 : tab2 = 23'b10000111111001011100111;
11'd1263 : tab2 = 23'b10000111101010010011101;
11'd1264 : tab2 = 23'b10000111011011001011010;
11'd1265 : tab2 = 23'b10000111001100000011111;
11'd1266 : tab2 = 23'b10000110111100111100110;
11'd1267 : tab2 = 23'b10000110101101110111001;
11'd1268 : tab2 = 23'b10000110011110110010011;
11'd1269 : tab2 = 23'b10000110001111101110000;
11'd1270 : tab2 = 23'b10000110000000101011001;
11'd1271 : tab2 = 23'b10000101110001101000100;
11'd1272 : tab2 = 23'b10000101100010100111001;
11'd1273 : tab2 = 23'b10000101010011100110101;
11'd1274 : tab2 = 23'b10000101000100100110110;
11'd1275 : tab2 = 23'b10000100110101100111110;
11'd1276 : tab2 = 23'b10000100100110101010000;
11'd1277 : tab2 = 23'b10000100010111101100110;
11'd1278 : tab2 = 23'b10000100001000110000100;
11'd1279 : tab2 = 23'b10000011111001110100111;
11'd1280 : tab2 = 23'b10000011101010111010011;
11'd1281 : tab2 = 23'b10000011011100000000111;
11'd1282 : tab2 = 23'b10000011001101001000001;
11'd1283 : tab2 = 23'b10000010111110001111110;
11'd1284 : tab2 = 23'b10000010101111011001000;
11'd1285 : tab2 = 23'b10000010100000100010011;
11'd1286 : tab2 = 23'b10000010010001101101011;
11'd1287 : tab2 = 23'b10000010000010111000100;
11'd1288 : tab2 = 23'b10000001110100000101000;
11'd1289 : tab2 = 23'b10000001100101010010000;
11'd1290 : tab2 = 23'b10000001010110100000010;
11'd1291 : tab2 = 23'b10000001000111101111000;
11'd1292 : tab2 = 23'b10000000111000111110110;
11'd1293 : tab2 = 23'b10000000101010001111011;
11'd1294 : tab2 = 23'b10000000011011100000101;
11'd1295 : tab2 = 23'b10000000001100110010101;
11'd1296 : tab2 = 23'b01111111111110000110000;
11'd1297 : tab2 = 23'b01111111101111011001111;
11'd1298 : tab2 = 23'b01111111100000101110101;
11'd1299 : tab2 = 23'b01111111010010000100010;
11'd1300 : tab2 = 23'b01111111000011011010111;
11'd1301 : tab2 = 23'b01111110110100110010000;
11'd1302 : tab2 = 23'b01111110100110001010000;
11'd1303 : tab2 = 23'b01111110010111100010111;
11'd1304 : tab2 = 23'b01111110001000111100110;
11'd1305 : tab2 = 23'b01111101111010010111100;
11'd1306 : tab2 = 23'b01111101101011110011000;
11'd1307 : tab2 = 23'b01111101011101001111100;
11'd1308 : tab2 = 23'b01111101001110101100010;
11'd1309 : tab2 = 23'b01111101000000001010100;
11'd1310 : tab2 = 23'b01111100110001101001000;
11'd1311 : tab2 = 23'b01111100100011001000110;
11'd1312 : tab2 = 23'b01111100010100101001011;
11'd1313 : tab2 = 23'b01111100000110001010101;
11'd1314 : tab2 = 23'b01111011110111101100101;
11'd1315 : tab2 = 23'b01111011101001001111101;
11'd1316 : tab2 = 23'b01111011011010110011100;
11'd1317 : tab2 = 23'b01111011001100011000001;
11'd1318 : tab2 = 23'b01111010111101111101001;
11'd1319 : tab2 = 23'b01111010101111100011101;
11'd1320 : tab2 = 23'b01111010100001001010110;
11'd1321 : tab2 = 23'b01111010010010110010110;
11'd1322 : tab2 = 23'b01111010000100011011010;
11'd1323 : tab2 = 23'b01111001110110000100101;
11'd1324 : tab2 = 23'b01111001100111101111010;
11'd1325 : tab2 = 23'b01111001011001011010001;
11'd1326 : tab2 = 23'b01111001001011000110001;
11'd1327 : tab2 = 23'b01111000111100110011000;
11'd1328 : tab2 = 23'b01111000101110100000111;
11'd1329 : tab2 = 23'b01111000100000001110111;
11'd1330 : tab2 = 23'b01111000010001111110001;
11'd1331 : tab2 = 23'b01111000000011101110010;
11'd1332 : tab2 = 23'b01110111110101011111000;
11'd1333 : tab2 = 23'b01110111100111010000101;
11'd1334 : tab2 = 23'b01110111011001000011000;
11'd1335 : tab2 = 23'b01110111001010110110011;
11'd1336 : tab2 = 23'b01110110111100101010100;
11'd1337 : tab2 = 23'b01110110101110011111000;
11'd1338 : tab2 = 23'b01110110100000010101000;
11'd1339 : tab2 = 23'b01110110010010001011100;
11'd1340 : tab2 = 23'b01110110000100000010111;
11'd1341 : tab2 = 23'b01110101110101111010111;
11'd1342 : tab2 = 23'b01110101100111110011101;
11'd1343 : tab2 = 23'b01110101011001101101011;
11'd1344 : tab2 = 23'b01110101001011100111111;
11'd1345 : tab2 = 23'b01110100111101100010110;
11'd1346 : tab2 = 23'b01110100101111011111000;
11'd1347 : tab2 = 23'b01110100100001011011111;
11'd1348 : tab2 = 23'b01110100010011011001101;
11'd1349 : tab2 = 23'b01110100000101011000000;
11'd1350 : tab2 = 23'b01110011110111010111001;
11'd1351 : tab2 = 23'b01110011101001010111001;
11'd1352 : tab2 = 23'b01110011011011011000001;
11'd1353 : tab2 = 23'b01110011001101011001111;
11'd1354 : tab2 = 23'b01110010111111011011111;
11'd1355 : tab2 = 23'b01110010110001011111011;
11'd1356 : tab2 = 23'b01110010100011100011001;
11'd1357 : tab2 = 23'b01110010010101101000000;
11'd1358 : tab2 = 23'b01110010000111101101100;
11'd1359 : tab2 = 23'b01110001111001110011111;
11'd1360 : tab2 = 23'b01110001101011111010110;
11'd1361 : tab2 = 23'b01110001011110000010111;
11'd1362 : tab2 = 23'b01110001010000001011100;
11'd1363 : tab2 = 23'b01110001000010010101000;
11'd1364 : tab2 = 23'b01110000110100011111000;
11'd1365 : tab2 = 23'b01110000100110101010010;
11'd1366 : tab2 = 23'b01110000011000110110000;
11'd1367 : tab2 = 23'b01110000001011000010011;
11'd1368 : tab2 = 23'b01101111111101001111111;
11'd1369 : tab2 = 23'b01101111101111011110010;
11'd1370 : tab2 = 23'b01101111100001101100110;
11'd1371 : tab2 = 23'b01101111010011111100101;
11'd1372 : tab2 = 23'b01101111000110001100111;
11'd1373 : tab2 = 23'b01101110111000011110000;
11'd1374 : tab2 = 23'b01101110101010110000001;
11'd1375 : tab2 = 23'b01101110011101000010101;
11'd1376 : tab2 = 23'b01101110001111010110011;
11'd1377 : tab2 = 23'b01101110000001101010011;
11'd1378 : tab2 = 23'b01101101110011111111100;
11'd1379 : tab2 = 23'b01101101100110010101100;
11'd1380 : tab2 = 23'b01101101011000101100001;
11'd1381 : tab2 = 23'b01101101001011000011100;
11'd1382 : tab2 = 23'b01101100111101011011001;
11'd1383 : tab2 = 23'b01101100101111110100010;
11'd1384 : tab2 = 23'b01101100100010001110000;
11'd1385 : tab2 = 23'b01101100010100101000100;
11'd1386 : tab2 = 23'b01101100000111000011100;
11'd1387 : tab2 = 23'b01101011111001011111011;
11'd1388 : tab2 = 23'b01101011101011111100001;
11'd1389 : tab2 = 23'b01101011011110011001010;
11'd1390 : tab2 = 23'b01101011010000110111101;
11'd1391 : tab2 = 23'b01101011000011010110011;
11'd1392 : tab2 = 23'b01101010110101110110010;
11'd1393 : tab2 = 23'b01101010101000010110101;
11'd1394 : tab2 = 23'b01101010011010110111111;
11'd1395 : tab2 = 23'b01101010001101011001101;
11'd1396 : tab2 = 23'b01101001111111111100101;
11'd1397 : tab2 = 23'b01101001110010011111110;
11'd1398 : tab2 = 23'b01101001100101000100001;
11'd1399 : tab2 = 23'b01101001010111101001000;
11'd1400 : tab2 = 23'b01101001001010001110101;
11'd1401 : tab2 = 23'b01101000111100110101000;
11'd1402 : tab2 = 23'b01101000101111011100011;
11'd1403 : tab2 = 23'b01101000100010000100010;
11'd1404 : tab2 = 23'b01101000010100101100110;
11'd1405 : tab2 = 23'b01101000000111010110011;
11'd1406 : tab2 = 23'b01100111111010000000101;
11'd1407 : tab2 = 23'b01100111101100101011101;
11'd1408 : tab2 = 23'b01100111011111010110111;
11'd1409 : tab2 = 23'b01100111010010000011010;
11'd1410 : tab2 = 23'b01100111000100110000100;
11'd1411 : tab2 = 23'b01100110110111011110010;
11'd1412 : tab2 = 23'b01100110101010001100111;
11'd1413 : tab2 = 23'b01100110011100111100011;
11'd1414 : tab2 = 23'b01100110001111101100000;
11'd1415 : tab2 = 23'b01100110000010011101001;
11'd1416 : tab2 = 23'b01100101110101001110100;
11'd1417 : tab2 = 23'b01100101101000000000110;
11'd1418 : tab2 = 23'b01100101011010110011110;
11'd1419 : tab2 = 23'b01100101001101100111101;
11'd1420 : tab2 = 23'b01100101000000011011110;
11'd1421 : tab2 = 23'b01100100110011010001010;
11'd1422 : tab2 = 23'b01100100100110000111000;
11'd1423 : tab2 = 23'b01100100011000111101101;
11'd1424 : tab2 = 23'b01100100001011110101001;
11'd1425 : tab2 = 23'b01100011111110101101001;
11'd1426 : tab2 = 23'b01100011110001100101111;
11'd1427 : tab2 = 23'b01100011100100011111010;
11'd1428 : tab2 = 23'b01100011010111011001110;
11'd1429 : tab2 = 23'b01100011001010010100100;
11'd1430 : tab2 = 23'b01100010111101010000010;
11'd1431 : tab2 = 23'b01100010110000001101000;
11'd1432 : tab2 = 23'b01100010100011001001111;
11'd1433 : tab2 = 23'b01100010010110000111111;
11'd1434 : tab2 = 23'b01100010001001000110001;
11'd1435 : tab2 = 23'b01100001111100000101101;
11'd1436 : tab2 = 23'b01100001101111000101110;
11'd1437 : tab2 = 23'b01100001100010000110010;
11'd1438 : tab2 = 23'b01100001010101000111111;
11'd1439 : tab2 = 23'b01100001001000001010000;
11'd1440 : tab2 = 23'b01100000111011001100111;
11'd1441 : tab2 = 23'b01100000101110010000011;
11'd1442 : tab2 = 23'b01100000100001010100111;
11'd1443 : tab2 = 23'b01100000010100011001110;
11'd1444 : tab2 = 23'b01100000000111011111011;
11'd1445 : tab2 = 23'b01011111111010100101111;
11'd1446 : tab2 = 23'b01011111101101101101001;
11'd1447 : tab2 = 23'b01011111100000110101000;
11'd1448 : tab2 = 23'b01011111010011111101101;
11'd1449 : tab2 = 23'b01011111000111000110110;
11'd1450 : tab2 = 23'b01011110111010010000110;
11'd1451 : tab2 = 23'b01011110101101011011101;
11'd1452 : tab2 = 23'b01011110100000100110101;
11'd1453 : tab2 = 23'b01011110010011110010110;
11'd1454 : tab2 = 23'b01011110000110111111110;
11'd1455 : tab2 = 23'b01011101111010001101010;
11'd1456 : tab2 = 23'b01011101101101011011000;
11'd1457 : tab2 = 23'b01011101100000101010001;
11'd1458 : tab2 = 23'b01011101010011111001110;
11'd1459 : tab2 = 23'b01011101000111001010000;
11'd1460 : tab2 = 23'b01011100111010011011000;
11'd1461 : tab2 = 23'b01011100101101101100100;
11'd1462 : tab2 = 23'b01011100100000111111001;
11'd1463 : tab2 = 23'b01011100010100010010000;
11'd1464 : tab2 = 23'b01011100000111100101110;
11'd1465 : tab2 = 23'b01011011111010111010010;
11'd1466 : tab2 = 23'b01011011101110001111100;
11'd1467 : tab2 = 23'b01011011100001100101011;
11'd1468 : tab2 = 23'b01011011010100111011110;
11'd1469 : tab2 = 23'b01011011001000010011001;
11'd1470 : tab2 = 23'b01011010111011101011001;
11'd1471 : tab2 = 23'b01011010101111000011011;
11'd1472 : tab2 = 23'b01011010100010011100111;
11'd1473 : tab2 = 23'b01011010010101110110110;
11'd1474 : tab2 = 23'b01011010001001010001011;
11'd1475 : tab2 = 23'b01011001111100101100111;
11'd1476 : tab2 = 23'b01011001110000001000111;
11'd1477 : tab2 = 23'b01011001100011100101101;
11'd1478 : tab2 = 23'b01011001010111000010111;
11'd1479 : tab2 = 23'b01011001001010100001000;
11'd1480 : tab2 = 23'b01011000111101111111111;
11'd1481 : tab2 = 23'b01011000110001011111000;
11'd1482 : tab2 = 23'b01011000100100111111010;
11'd1483 : tab2 = 23'b01011000011000100000000;
11'd1484 : tab2 = 23'b01011000001100000001010;
11'd1485 : tab2 = 23'b01010111111111100011101;
11'd1486 : tab2 = 23'b01010111110011000110100;
11'd1487 : tab2 = 23'b01010111100110101001111;
11'd1488 : tab2 = 23'b01010111011010001110011;
11'd1489 : tab2 = 23'b01010111001101110010111;
11'd1490 : tab2 = 23'b01010111000001011000101;
11'd1491 : tab2 = 23'b01010110110100111110101;
11'd1492 : tab2 = 23'b01010110101000100101100;
11'd1493 : tab2 = 23'b01010110011100001101001;
11'd1494 : tab2 = 23'b01010110001111110101101;
11'd1495 : tab2 = 23'b01010110000011011110010;
11'd1496 : tab2 = 23'b01010101110111001000000;
11'd1497 : tab2 = 23'b01010101101010110010000;
11'd1498 : tab2 = 23'b01010101011110011101000;
11'd1499 : tab2 = 23'b01010101010010001000101;
11'd1500 : tab2 = 23'b01010101000101110100110;
11'd1501 : tab2 = 23'b01010100111001100001111;
11'd1502 : tab2 = 23'b01010100101101001111100;
11'd1503 : tab2 = 23'b01010100100000111101100;
11'd1504 : tab2 = 23'b01010100010100101100100;
11'd1505 : tab2 = 23'b01010100001000011100000;
11'd1506 : tab2 = 23'b01010011111100001100000;
11'd1507 : tab2 = 23'b01010011101111111101000;
11'd1508 : tab2 = 23'b01010011100011101110101;
11'd1509 : tab2 = 23'b01010011010111100000110;
11'd1510 : tab2 = 23'b01010011001011010011011;
11'd1511 : tab2 = 23'b01010010111111000111001;
11'd1512 : tab2 = 23'b01010010110010111011010;
11'd1513 : tab2 = 23'b01010010100110110000010;
11'd1514 : tab2 = 23'b01010010011010100101110;
11'd1515 : tab2 = 23'b01010010001110011011100;
11'd1516 : tab2 = 23'b01010010000010010010101;
11'd1517 : tab2 = 23'b01010001110110001001111;
11'd1518 : tab2 = 23'b01010001101010000010000;
11'd1519 : tab2 = 23'b01010001011101111010111;
11'd1520 : tab2 = 23'b01010001010001110100011;
11'd1521 : tab2 = 23'b01010001000101101110010;
11'd1522 : tab2 = 23'b01010000111001101001010;
11'd1523 : tab2 = 23'b01010000101101100100001;
11'd1524 : tab2 = 23'b01010000100001100000011;
11'd1525 : tab2 = 23'b01010000010101011100111;
11'd1526 : tab2 = 23'b01010000001001011010001;
11'd1527 : tab2 = 23'b01001111111101011000010;
11'd1528 : tab2 = 23'b01001111110001010110110;
11'd1529 : tab2 = 23'b01001111100101010110001;
11'd1530 : tab2 = 23'b01001111011001010110000;
11'd1531 : tab2 = 23'b01001111001101010110101;
11'd1532 : tab2 = 23'b01001111000001010111100;
11'd1533 : tab2 = 23'b01001110110101011001100;
11'd1534 : tab2 = 23'b01001110101001011011111;
11'd1535 : tab2 = 23'b01001110011101011110110;
11'd1536 : tab2 = 23'b01001110010001100010110;
11'd1537 : tab2 = 23'b01001110000101100111000;
11'd1538 : tab2 = 23'b01001101111001101100000;
11'd1539 : tab2 = 23'b01001101101101110001110;
11'd1540 : tab2 = 23'b01001101100001111000001;
11'd1541 : tab2 = 23'b01001101010101111111001;
11'd1542 : tab2 = 23'b01001101001010000110110;
11'd1543 : tab2 = 23'b01001100111110001110110;
11'd1544 : tab2 = 23'b01001100110010010111101;
11'd1545 : tab2 = 23'b01001100100110100000111;
11'd1546 : tab2 = 23'b01001100011010101011000;
11'd1547 : tab2 = 23'b01001100001110110101111;
11'd1548 : tab2 = 23'b01001100000011000001000;
11'd1549 : tab2 = 23'b01001011110111001101010;
11'd1550 : tab2 = 23'b01001011101011011001101;
11'd1551 : tab2 = 23'b01001011011111100111000;
11'd1552 : tab2 = 23'b01001011010011110101000;
11'd1553 : tab2 = 23'b01001011001000000011011;
11'd1554 : tab2 = 23'b01001010111100010010011;
11'd1555 : tab2 = 23'b01001010110000100010010;
11'd1556 : tab2 = 23'b01001010100100110010110;
11'd1557 : tab2 = 23'b01001010011001000011110;
11'd1558 : tab2 = 23'b01001010001101010101010;
11'd1559 : tab2 = 23'b01001010000001100111110;
11'd1560 : tab2 = 23'b01001001110101111010100;
11'd1561 : tab2 = 23'b01001001101010001110000;
11'd1562 : tab2 = 23'b01001001011110100010010;
11'd1563 : tab2 = 23'b01001001010010110110110;
11'd1564 : tab2 = 23'b01001001000111001100010;
11'd1565 : tab2 = 23'b01001000111011100010000;
11'd1566 : tab2 = 23'b01001000101111111000111;
11'd1567 : tab2 = 23'b01001000100100010000001;
11'd1568 : tab2 = 23'b01001000011000101000000;
11'd1569 : tab2 = 23'b01001000001101000000010;
11'd1570 : tab2 = 23'b01001000000001011001100;
11'd1571 : tab2 = 23'b01000111110101110011001;
11'd1572 : tab2 = 23'b01000111101010001101011;
11'd1573 : tab2 = 23'b01000111011110101000100;
11'd1574 : tab2 = 23'b01000111010011000011110;
11'd1575 : tab2 = 23'b01000111000111100000001;
11'd1576 : tab2 = 23'b01000110111011111100101;
11'd1577 : tab2 = 23'b01000110110000011010010;
11'd1578 : tab2 = 23'b01000110100100111000000;
11'd1579 : tab2 = 23'b01000110011001010110101;
11'd1580 : tab2 = 23'b01000110001101110101111;
11'd1581 : tab2 = 23'b01000110000010010101110;
11'd1582 : tab2 = 23'b01000101110110110110010;
11'd1583 : tab2 = 23'b01000101101011010111011;
11'd1584 : tab2 = 23'b01000101011111111000101;
11'd1585 : tab2 = 23'b01000101010100011011000;
11'd1586 : tab2 = 23'b01000101001000111110000;
11'd1587 : tab2 = 23'b01000100111101100001101;
11'd1588 : tab2 = 23'b01000100110010000101011;
11'd1589 : tab2 = 23'b01000100100110101010001;
11'd1590 : tab2 = 23'b01000100011011001111010;
11'd1591 : tab2 = 23'b01000100001111110101010;
11'd1592 : tab2 = 23'b01000100000100011011110;
11'd1593 : tab2 = 23'b01000011111001000010111;
11'd1594 : tab2 = 23'b01000011101101101010011;
11'd1595 : tab2 = 23'b01000011100010010010111;
11'd1596 : tab2 = 23'b01000011010110111011101;
11'd1597 : tab2 = 23'b01000011001011100101001;
11'd1598 : tab2 = 23'b01000011000000001111001;
11'd1599 : tab2 = 23'b01000010110100111001111;
11'd1600 : tab2 = 23'b01000010101001100101001;
11'd1601 : tab2 = 23'b01000010011110010001001;
11'd1602 : tab2 = 23'b01000010010010111101010;
11'd1603 : tab2 = 23'b01000010000111101010010;
11'd1604 : tab2 = 23'b01000001111100010111111;
11'd1605 : tab2 = 23'b01000001110001000110011;
11'd1606 : tab2 = 23'b01000001100101110101000;
11'd1607 : tab2 = 23'b01000001011010100100100;
11'd1608 : tab2 = 23'b01000001001111010100101;
11'd1609 : tab2 = 23'b01000001000100000101000;
11'd1610 : tab2 = 23'b01000000111000110110001;
11'd1611 : tab2 = 23'b01000000101101101000000;
11'd1612 : tab2 = 23'b01000000100010011010011;
11'd1613 : tab2 = 23'b01000000010111001101010;
11'd1614 : tab2 = 23'b01000000001100000000110;
11'd1615 : tab2 = 23'b01000000000000110100111;
11'd1616 : tab2 = 23'b00111111110101101001101;
11'd1617 : tab2 = 23'b00111111101010011110110;
11'd1618 : tab2 = 23'b00111111011111010100110;
11'd1619 : tab2 = 23'b00111111010100001011010;
11'd1620 : tab2 = 23'b00111111001001000010010;
11'd1621 : tab2 = 23'b00111110111101111001110;
11'd1622 : tab2 = 23'b00111110110010110010010;
11'd1623 : tab2 = 23'b00111110100111101011000;
11'd1624 : tab2 = 23'b00111110011100100100011;
11'd1625 : tab2 = 23'b00111110010001011110010;
11'd1626 : tab2 = 23'b00111110000110011000110;
11'd1627 : tab2 = 23'b00111101111011010100001;
11'd1628 : tab2 = 23'b00111101110000001111100;
11'd1629 : tab2 = 23'b00111101100101001011110;
11'd1630 : tab2 = 23'b00111101011010001000111;
11'd1631 : tab2 = 23'b00111101001111000110000;
11'd1632 : tab2 = 23'b00111101000100000100010;
11'd1633 : tab2 = 23'b00111100111001000010110;
11'd1634 : tab2 = 23'b00111100101110000010001;
11'd1635 : tab2 = 23'b00111100100011000001100;
11'd1636 : tab2 = 23'b00111100011000000001110;
11'd1637 : tab2 = 23'b00111100001101000010110;
11'd1638 : tab2 = 23'b00111100000010000100001;
11'd1639 : tab2 = 23'b00111011110111000110010;
11'd1640 : tab2 = 23'b00111011101100001000111;
11'd1641 : tab2 = 23'b00111011100001001011110;
11'd1642 : tab2 = 23'b00111011010110001111101;
11'd1643 : tab2 = 23'b00111011001011010011111;
11'd1644 : tab2 = 23'b00111011000000011000110;
11'd1645 : tab2 = 23'b00111010110101011110010;
11'd1646 : tab2 = 23'b00111010101010100100010;
11'd1647 : tab2 = 23'b00111010011111101010110;
11'd1648 : tab2 = 23'b00111010010100110001111;
11'd1649 : tab2 = 23'b00111010001001111001100;
11'd1650 : tab2 = 23'b00111001111111000001110;
11'd1651 : tab2 = 23'b00111001110100001010101;
11'd1652 : tab2 = 23'b00111001101001010100010;
11'd1653 : tab2 = 23'b00111001011110011110000;
11'd1654 : tab2 = 23'b00111001010011101000100;
11'd1655 : tab2 = 23'b00111001001000110011100;
11'd1656 : tab2 = 23'b00111000111101111111010;
11'd1657 : tab2 = 23'b00111000110011001011100;
11'd1658 : tab2 = 23'b00111000101000011000001;
11'd1659 : tab2 = 23'b00111000011101100101011;
11'd1660 : tab2 = 23'b00111000010010110011100;
11'd1661 : tab2 = 23'b00111000001000000001111;
11'd1662 : tab2 = 23'b00110111111101010000111;
11'd1663 : tab2 = 23'b00110111110010100000001;
11'd1664 : tab2 = 23'b00110111100111110000011;
11'd1665 : tab2 = 23'b00110111011101000000111;
11'd1666 : tab2 = 23'b00110111010010010010011;
11'd1667 : tab2 = 23'b00110111000111100100000;
11'd1668 : tab2 = 23'b00110110111100110110011;
11'd1669 : tab2 = 23'b00110110110010001001010;
11'd1670 : tab2 = 23'b00110110100111011100101;
11'd1671 : tab2 = 23'b00110110011100110000011;
11'd1672 : tab2 = 23'b00110110010010000101001;
11'd1673 : tab2 = 23'b00110110000111011010001;
11'd1674 : tab2 = 23'b00110101111100101111110;
11'd1675 : tab2 = 23'b00110101110010000110000;
11'd1676 : tab2 = 23'b00110101100111011100111;
11'd1677 : tab2 = 23'b00110101011100110100010;
11'd1678 : tab2 = 23'b00110101010010001011110;
11'd1679 : tab2 = 23'b00110101000111100100010;
11'd1680 : tab2 = 23'b00110100111100111101000;
11'd1681 : tab2 = 23'b00110100110010010110110;
11'd1682 : tab2 = 23'b00110100100111110000101;
11'd1683 : tab2 = 23'b00110100011101001011010;
11'd1684 : tab2 = 23'b00110100010010100110001;
11'd1685 : tab2 = 23'b00110100001000000001111;
11'd1686 : tab2 = 23'b00110011111101011101111;
11'd1687 : tab2 = 23'b00110011110010111010111;
11'd1688 : tab2 = 23'b00110011101000011000001;
11'd1689 : tab2 = 23'b00110011011101110110000;
11'd1690 : tab2 = 23'b00110011010011010100001;
11'd1691 : tab2 = 23'b00110011001000110011000;
11'd1692 : tab2 = 23'b00110010111110010010100;
11'd1693 : tab2 = 23'b00110010110011110010100;
11'd1694 : tab2 = 23'b00110010101001010011010;
11'd1695 : tab2 = 23'b00110010011110110011111;
11'd1696 : tab2 = 23'b00110010010100010101111;
11'd1697 : tab2 = 23'b00110010001001110111111;
11'd1698 : tab2 = 23'b00110001111111011010100;
11'd1699 : tab2 = 23'b00110001110100111101110;
11'd1700 : tab2 = 23'b00110001101010100001100;
11'd1701 : tab2 = 23'b00110001100000000101101;
11'd1702 : tab2 = 23'b00110001010101101010100;
11'd1703 : tab2 = 23'b00110001001011001111111;
11'd1704 : tab2 = 23'b00110001000000110101101;
11'd1705 : tab2 = 23'b00110000110110011100010;
11'd1706 : tab2 = 23'b00110000101100000011001;
11'd1707 : tab2 = 23'b00110000100001101010011;
11'd1708 : tab2 = 23'b00110000010111010010100;
11'd1709 : tab2 = 23'b00110000001100111010110;
11'd1710 : tab2 = 23'b00110000000010100100001;
11'd1711 : tab2 = 23'b00101111111000001101101;
11'd1712 : tab2 = 23'b00101111101101110111110;
11'd1713 : tab2 = 23'b00101111100011100010100;
11'd1714 : tab2 = 23'b00101111011001001101101;
11'd1715 : tab2 = 23'b00101111001110111001001;
11'd1716 : tab2 = 23'b00101111000100100101011;
11'd1717 : tab2 = 23'b00101110111010010010011;
11'd1718 : tab2 = 23'b00101110101111111111010;
11'd1719 : tab2 = 23'b00101110100101101101010;
11'd1720 : tab2 = 23'b00101110011011011011110;
11'd1721 : tab2 = 23'b00101110010001001010011;
11'd1722 : tab2 = 23'b00101110000110111001111;
11'd1723 : tab2 = 23'b00101101111100101001100;
11'd1724 : tab2 = 23'b00101101110010011010001;
11'd1725 : tab2 = 23'b00101101101000001011000;
11'd1726 : tab2 = 23'b00101101011101111100100;
11'd1727 : tab2 = 23'b00101101010011101110010;
11'd1728 : tab2 = 23'b00101101001001100000110;
11'd1729 : tab2 = 23'b00101100111111010011111;
11'd1730 : tab2 = 23'b00101100110101000111100;
11'd1731 : tab2 = 23'b00101100101010111011010;
11'd1732 : tab2 = 23'b00101100100000110000000;
11'd1733 : tab2 = 23'b00101100010110100101010;
11'd1734 : tab2 = 23'b00101100001100011010100;
11'd1735 : tab2 = 23'b00101100000010010000111;
11'd1736 : tab2 = 23'b00101011111000000111100;
11'd1737 : tab2 = 23'b00101011101101111110110;
11'd1738 : tab2 = 23'b00101011100011110110001;
11'd1739 : tab2 = 23'b00101011011001101110010;
11'd1740 : tab2 = 23'b00101011001111100111000;
11'd1741 : tab2 = 23'b00101011000101100000011;
11'd1742 : tab2 = 23'b00101010111011011001110;
11'd1743 : tab2 = 23'b00101010110001010100010;
11'd1744 : tab2 = 23'b00101010100111001110111;
11'd1745 : tab2 = 23'b00101010011101001010001;
11'd1746 : tab2 = 23'b00101010010011000101111;
11'd1747 : tab2 = 23'b00101010001001000010011;
11'd1748 : tab2 = 23'b00101001111110111110110;
11'd1749 : tab2 = 23'b00101001110100111100010;
11'd1750 : tab2 = 23'b00101001101010111010001;
11'd1751 : tab2 = 23'b00101001100000111000010;
11'd1752 : tab2 = 23'b00101001010110110111000;
11'd1753 : tab2 = 23'b00101001001100110110101;
11'd1754 : tab2 = 23'b00101001000010110110001;
11'd1755 : tab2 = 23'b00101000111000110110011;
11'd1756 : tab2 = 23'b00101000101110110111010;
11'd1757 : tab2 = 23'b00101000100100111000101;
11'd1758 : tab2 = 23'b00101000011010111010010;
11'd1759 : tab2 = 23'b00101000010000111100110;
11'd1760 : tab2 = 23'b00101000000110111111011;
11'd1761 : tab2 = 23'b00100111111101000010110;
11'd1762 : tab2 = 23'b00100111110011000110101;
11'd1763 : tab2 = 23'b00100111101001001011001;
11'd1764 : tab2 = 23'b00100111011111001111101;
11'd1765 : tab2 = 23'b00100111010101010101010;
11'd1766 : tab2 = 23'b00100111001011011011001;
11'd1767 : tab2 = 23'b00100111000001100001011;
11'd1768 : tab2 = 23'b00100110110111101000001;
11'd1769 : tab2 = 23'b00100110101101101111010;
11'd1770 : tab2 = 23'b00100110100011110111011;
11'd1771 : tab2 = 23'b00100110011001111111101;
11'd1772 : tab2 = 23'b00100110010000001000011;
11'd1773 : tab2 = 23'b00100110000110010001110;
11'd1774 : tab2 = 23'b00100101111100011011101;
11'd1775 : tab2 = 23'b00100101110010100101111;
11'd1776 : tab2 = 23'b00100101101000110000101;
11'd1777 : tab2 = 23'b00100101011110111011110;
11'd1778 : tab2 = 23'b00100101010101000111101;
11'd1779 : tab2 = 23'b00100101001011010100001;
11'd1780 : tab2 = 23'b00100101000001100000100;
11'd1781 : tab2 = 23'b00100100110111101110000;
11'd1782 : tab2 = 23'b00100100101101111011100;
11'd1783 : tab2 = 23'b00100100100100001001110;
11'd1784 : tab2 = 23'b00100100011010011000110;
11'd1785 : tab2 = 23'b00100100010000100111111;
11'd1786 : tab2 = 23'b00100100000110110111100;
11'd1787 : tab2 = 23'b00100011111101000111110;
11'd1788 : tab2 = 23'b00100011110011011000011;
11'd1789 : tab2 = 23'b00100011101001101001100;
11'd1790 : tab2 = 23'b00100011011111111011010;
11'd1791 : tab2 = 23'b00100011010110001101010;
11'd1792 : tab2 = 23'b00100011001100100000000;
11'd1793 : tab2 = 23'b00100011000010110011000;
11'd1794 : tab2 = 23'b00100010111001000110111;
11'd1795 : tab2 = 23'b00100010101111011010100;
11'd1796 : tab2 = 23'b00100010100101101111011;
11'd1797 : tab2 = 23'b00100010011100000100100;
11'd1798 : tab2 = 23'b00100010010010011001110;
11'd1799 : tab2 = 23'b00100010001000101111111;
11'd1800 : tab2 = 23'b00100001111111000110010;
11'd1801 : tab2 = 23'b00100001110101011101011;
11'd1802 : tab2 = 23'b00100001101011110100100;
11'd1803 : tab2 = 23'b00100001100010001100110;
11'd1804 : tab2 = 23'b00100001011000100101000;
11'd1805 : tab2 = 23'b00100001001110111110000;
11'd1806 : tab2 = 23'b00100001000101010111100;
11'd1807 : tab2 = 23'b00100000111011110001001;
11'd1808 : tab2 = 23'b00100000110010001011101;
11'd1809 : tab2 = 23'b00100000101000100110011;
11'd1810 : tab2 = 23'b00100000011111000001110;
11'd1811 : tab2 = 23'b00100000010101011101011;
11'd1812 : tab2 = 23'b00100000001011111001101;
11'd1813 : tab2 = 23'b00100000000010010110010;
11'd1814 : tab2 = 23'b00011111111000110011101;
11'd1815 : tab2 = 23'b00011111101111010001001;
11'd1816 : tab2 = 23'b00011111100101101111011;
11'd1817 : tab2 = 23'b00011111011100001110000;
11'd1818 : tab2 = 23'b00011111010010101101000;
11'd1819 : tab2 = 23'b00011111001001001100100;
11'd1820 : tab2 = 23'b00011110111111101100011;
11'd1821 : tab2 = 23'b00011110110110001101000;
11'd1822 : tab2 = 23'b00011110101100101101110;
11'd1823 : tab2 = 23'b00011110100011001111100;
11'd1824 : tab2 = 23'b00011110011001110001010;
11'd1825 : tab2 = 23'b00011110010000010011111;
11'd1826 : tab2 = 23'b00011110000110110110100;
11'd1827 : tab2 = 23'b00011101111101011001111;
11'd1828 : tab2 = 23'b00011101110011111101110;
11'd1829 : tab2 = 23'b00011101101010100001101;
11'd1830 : tab2 = 23'b00011101100001000110100;
11'd1831 : tab2 = 23'b00011101010111101011101;
11'd1832 : tab2 = 23'b00011101001110010001011;
11'd1833 : tab2 = 23'b00011101000100110111100;
11'd1834 : tab2 = 23'b00011100111011011101111;
11'd1835 : tab2 = 23'b00011100110010000101001;
11'd1836 : tab2 = 23'b00011100101000101100100;
11'd1837 : tab2 = 23'b00011100011111010100101;
11'd1838 : tab2 = 23'b00011100010101111100111;
11'd1839 : tab2 = 23'b00011100001100100101110;
11'd1840 : tab2 = 23'b00011100000011001111001;
11'd1841 : tab2 = 23'b00011011111001111001001;
11'd1842 : tab2 = 23'b00011011110000100011011;
11'd1843 : tab2 = 23'b00011011100111001110010;
11'd1844 : tab2 = 23'b00011011011101111001010;
11'd1845 : tab2 = 23'b00011011010100100100111;
11'd1846 : tab2 = 23'b00011011001011010001000;
11'd1847 : tab2 = 23'b00011011000001111101100;
11'd1848 : tab2 = 23'b00011010111000101010110;
11'd1849 : tab2 = 23'b00011010101111011000001;
11'd1850 : tab2 = 23'b00011010100110000110001;
11'd1851 : tab2 = 23'b00011010011100110100101;
11'd1852 : tab2 = 23'b00011010010011100011010;
11'd1853 : tab2 = 23'b00011010001010010010100;
11'd1854 : tab2 = 23'b00011010000001000010100;
11'd1855 : tab2 = 23'b00011001110111110010101;
11'd1856 : tab2 = 23'b00011001101110100011011;
11'd1857 : tab2 = 23'b00011001100101010100101;
11'd1858 : tab2 = 23'b00011001011100000101111;
11'd1859 : tab2 = 23'b00011001010010111000010;
11'd1860 : tab2 = 23'b00011001001001101010101;
11'd1861 : tab2 = 23'b00011001000000011101100;
11'd1862 : tab2 = 23'b00011000110111010001000;
11'd1863 : tab2 = 23'b00011000101110000101000;
11'd1864 : tab2 = 23'b00011000100100111001000;
11'd1865 : tab2 = 23'b00011000011011101101111;
11'd1866 : tab2 = 23'b00011000010010100011000;
11'd1867 : tab2 = 23'b00011000001001011000111;
11'd1868 : tab2 = 23'b00011000000000001110111;
11'd1869 : tab2 = 23'b00010111110111000101100;
11'd1870 : tab2 = 23'b00010111101101111100101;
11'd1871 : tab2 = 23'b00010111100100110011111;
11'd1872 : tab2 = 23'b00010111011011101011110;
11'd1873 : tab2 = 23'b00010111010010100100000;
11'd1874 : tab2 = 23'b00010111001001011101000;
11'd1875 : tab2 = 23'b00010111000000010101111;
11'd1876 : tab2 = 23'b00010110110111001111110;
11'd1877 : tab2 = 23'b00010110101110001001101;
11'd1878 : tab2 = 23'b00010110100101000100100;
11'd1879 : tab2 = 23'b00010110011011111111100;
11'd1880 : tab2 = 23'b00010110010010111011000;
11'd1881 : tab2 = 23'b00010110001001110110111;
11'd1882 : tab2 = 23'b00010110000000110011001;
11'd1883 : tab2 = 23'b00010101110111101111110;
11'd1884 : tab2 = 23'b00010101101110101101001;
11'd1885 : tab2 = 23'b00010101100101101010111;
11'd1886 : tab2 = 23'b00010101011100101000110;
11'd1887 : tab2 = 23'b00010101010011100111100;
11'd1888 : tab2 = 23'b00010101001010100110100;
11'd1889 : tab2 = 23'b00010101000001100101111;
11'd1890 : tab2 = 23'b00010100111000100101111;
11'd1891 : tab2 = 23'b00010100101111100110000;
11'd1892 : tab2 = 23'b00010100100110100110111;
11'd1893 : tab2 = 23'b00010100011101101000001;
11'd1894 : tab2 = 23'b00010100010100101001100;
11'd1895 : tab2 = 23'b00010100001011101011101;
11'd1896 : tab2 = 23'b00010100000010101110001;
11'd1897 : tab2 = 23'b00010011111001110001010;
11'd1898 : tab2 = 23'b00010011110000110100100;
11'd1899 : tab2 = 23'b00010011100111111000011;
11'd1900 : tab2 = 23'b00010011011110111100100;
11'd1901 : tab2 = 23'b00010011010110000001010;
11'd1902 : tab2 = 23'b00010011001101000110011;
11'd1903 : tab2 = 23'b00010011000100001011110;
11'd1904 : tab2 = 23'b00010010111011010001101;
11'd1905 : tab2 = 23'b00010010110010011000010;
11'd1906 : tab2 = 23'b00010010101001011111000;
11'd1907 : tab2 = 23'b00010010100000100110010;
11'd1908 : tab2 = 23'b00010010010111101110000;
11'd1909 : tab2 = 23'b00010010001110110110010;
11'd1910 : tab2 = 23'b00010010000101111110101;
11'd1911 : tab2 = 23'b00010001111101000111110;
11'd1912 : tab2 = 23'b00010001110100010001001;
11'd1913 : tab2 = 23'b00010001101011011010110;
11'd1914 : tab2 = 23'b00010001100010100101010;
11'd1915 : tab2 = 23'b00010001011001101111111;
11'd1916 : tab2 = 23'b00010001010000111011001;
11'd1917 : tab2 = 23'b00010001001000000110101;
11'd1918 : tab2 = 23'b00010000111111010010110;
11'd1919 : tab2 = 23'b00010000110110011111000;
11'd1920 : tab2 = 23'b00010000101101101011111;
11'd1921 : tab2 = 23'b00010000100100111000111;
11'd1922 : tab2 = 23'b00010000011100000110101;
11'd1923 : tab2 = 23'b00010000010011010101000;
11'd1924 : tab2 = 23'b00010000001010100011100;
11'd1925 : tab2 = 23'b00010000000001110010011;
11'd1926 : tab2 = 23'b00001111111001000001101;
11'd1927 : tab2 = 23'b00001111110000010001011;
11'd1928 : tab2 = 23'b00001111100111100001110;
11'd1929 : tab2 = 23'b00001111011110110010010;
11'd1930 : tab2 = 23'b00001111010110000011101;
11'd1931 : tab2 = 23'b00001111001101010101001;
11'd1932 : tab2 = 23'b00001111000100100110111;
11'd1933 : tab2 = 23'b00001110111011111001010;
11'd1934 : tab2 = 23'b00001110110011001100000;
11'd1935 : tab2 = 23'b00001110101010011111011;
11'd1936 : tab2 = 23'b00001110100001110010101;
11'd1937 : tab2 = 23'b00001110011001000110100;
11'd1938 : tab2 = 23'b00001110010000011011001;
11'd1939 : tab2 = 23'b00001110000111101111111;
11'd1940 : tab2 = 23'b00001101111111000101010;
11'd1941 : tab2 = 23'b00001101110110011011000;
11'd1942 : tab2 = 23'b00001101101101110000111;
11'd1943 : tab2 = 23'b00001101100101000111110;
11'd1944 : tab2 = 23'b00001101011100011110101;
11'd1945 : tab2 = 23'b00001101010011110101110;
11'd1946 : tab2 = 23'b00001101001011001101100;
11'd1947 : tab2 = 23'b00001101000010100101111;
11'd1948 : tab2 = 23'b00001100111001111110100;
11'd1949 : tab2 = 23'b00001100110001010111011;
11'd1950 : tab2 = 23'b00001100101000110001000;
11'd1951 : tab2 = 23'b00001100100000001010110;
11'd1952 : tab2 = 23'b00001100010111100101000;
11'd1953 : tab2 = 23'b00001100001110111111101;
11'd1954 : tab2 = 23'b00001100000110011010110;
11'd1955 : tab2 = 23'b00001011111101110110010;
11'd1956 : tab2 = 23'b00001011110101010010000;
11'd1957 : tab2 = 23'b00001011101100101110010;
11'd1958 : tab2 = 23'b00001011100100001011000;
11'd1959 : tab2 = 23'b00001011011011101000001;
11'd1960 : tab2 = 23'b00001011010011000101101;
11'd1961 : tab2 = 23'b00001011001010100011100;
11'd1962 : tab2 = 23'b00001011000010000010001;
11'd1963 : tab2 = 23'b00001010111001100000110;
11'd1964 : tab2 = 23'b00001010110000111111111;
11'd1965 : tab2 = 23'b00001010101000011111101;
11'd1966 : tab2 = 23'b00001010011111111111011;
11'd1967 : tab2 = 23'b00001010010111011111111;
11'd1968 : tab2 = 23'b00001010001111000000100;
11'd1969 : tab2 = 23'b00001010000110100001111;
11'd1970 : tab2 = 23'b00001001111110000011100;
11'd1971 : tab2 = 23'b00001001110101100101011;
11'd1972 : tab2 = 23'b00001001101101000111110;
11'd1973 : tab2 = 23'b00001001100100101010101;
11'd1974 : tab2 = 23'b00001001011100001101101;
11'd1975 : tab2 = 23'b00001001010011110001100;
11'd1976 : tab2 = 23'b00001001001011010101100;
11'd1977 : tab2 = 23'b00001001000010111001111;
11'd1978 : tab2 = 23'b00001000111010011110111;
11'd1979 : tab2 = 23'b00001000110010000011111;
11'd1980 : tab2 = 23'b00001000101001101001011;
11'd1981 : tab2 = 23'b00001000100001001111101;
11'd1982 : tab2 = 23'b00001000011000110101111;
11'd1983 : tab2 = 23'b00001000010000011100111;
11'd1984 : tab2 = 23'b00001000001000000100000;
11'd1985 : tab2 = 23'b00000111111111101011110;
11'd1986 : tab2 = 23'b00000111110111010011101;
11'd1987 : tab2 = 23'b00000111101110111100001;
11'd1988 : tab2 = 23'b00000111100110100100111;
11'd1989 : tab2 = 23'b00000111011110001110001;
11'd1990 : tab2 = 23'b00000111010101110111111;
11'd1991 : tab2 = 23'b00000111001101100001101;
11'd1992 : tab2 = 23'b00000111000101001100011;
11'd1993 : tab2 = 23'b00000110111100110111001;
11'd1994 : tab2 = 23'b00000110110100100010001;
11'd1995 : tab2 = 23'b00000110101100001101110;
11'd1996 : tab2 = 23'b00000110100011111001110;
11'd1997 : tab2 = 23'b00000110011011100110011;
11'd1998 : tab2 = 23'b00000110010011010010111;
11'd1999 : tab2 = 23'b00000110001011000000000;
11'd2000 : tab2 = 23'b00000110000010101101111;
11'd2001 : tab2 = 23'b00000101111010011011110;
11'd2002 : tab2 = 23'b00000101110010001010001;
11'd2003 : tab2 = 23'b00000101101001111001000;
11'd2004 : tab2 = 23'b00000101100001101000001;
11'd2005 : tab2 = 23'b00000101011001010111100;
11'd2006 : tab2 = 23'b00000101010001000111011;
11'd2007 : tab2 = 23'b00000101001000110111101;
11'd2008 : tab2 = 23'b00000101000000101000011;
11'd2009 : tab2 = 23'b00000100111000011001011;
11'd2010 : tab2 = 23'b00000100110000001011000;
11'd2011 : tab2 = 23'b00000100100111111100110;
11'd2012 : tab2 = 23'b00000100011111101111001;
11'd2013 : tab2 = 23'b00000100010111100001101;
11'd2014 : tab2 = 23'b00000100001111010100110;
11'd2015 : tab2 = 23'b00000100000111001000011;
11'd2016 : tab2 = 23'b00000011111110111100000;
11'd2017 : tab2 = 23'b00000011110110110000010;
11'd2018 : tab2 = 23'b00000011101110100100101;
11'd2019 : tab2 = 23'b00000011100110011001110;
11'd2020 : tab2 = 23'b00000011011110001111001;
11'd2021 : tab2 = 23'b00000011010110000101000;
11'd2022 : tab2 = 23'b00000011001101111011001;
11'd2023 : tab2 = 23'b00000011000101110001100;
11'd2024 : tab2 = 23'b00000010111101101000011;
11'd2025 : tab2 = 23'b00000010110101011111110;
11'd2026 : tab2 = 23'b00000010101101010111010;
11'd2027 : tab2 = 23'b00000010100101001111100;
11'd2028 : tab2 = 23'b00000010011101001000000;
11'd2029 : tab2 = 23'b00000010010101000000101;
11'd2030 : tab2 = 23'b00000010001100111001110;
11'd2031 : tab2 = 23'b00000010000100110011011;
11'd2032 : tab2 = 23'b00000001111100101101011;
11'd2033 : tab2 = 23'b00000001110100100111110;
11'd2034 : tab2 = 23'b00000001101100100010100;
11'd2035 : tab2 = 23'b00000001100100011101101;
11'd2036 : tab2 = 23'b00000001011100011000110;
11'd2037 : tab2 = 23'b00000001010100010100111;
11'd2038 : tab2 = 23'b00000001001100010001001;
11'd2039 : tab2 = 23'b00000001000100001101110;
11'd2040 : tab2 = 23'b00000000111100001010100;
11'd2041 : tab2 = 23'b00000000110100001000001;
11'd2042 : tab2 = 23'b00000000101100000101111;
11'd2043 : tab2 = 23'b00000000100100000100000;
11'd2044 : tab2 = 23'b00000000011100000010010;
11'd2045 : tab2 = 23'b00000000010100000001011;
11'd2046 : tab2 = 23'b00000000001100000000101;
11'd2047 : tab2 = 23'b00000000000100000000010;
endcase
  end
  endfunction

  wire [0:0] swire;
  wire [7:0] ewire;
  wire [22:0] m;

  assign swire = x[31];
  assign ewire = x[30:23];
  assign m = x[22:0];

  wire [23:0] mawire;

  wire [22:0] x0wire;
  
  assign x0wire = tab(m[22:12]);

  assign mawire = (ewire == 8'b0) ? {1'b0,m[22:0]} : {1'b1,m[22:0]};
  
  wire [22:0] x2wire;


  reg [22:0] x0reg;
  reg [23:0] mareg;
  reg [22:0] x2reg;
  reg [7:0] ereg;
  reg sreg;
  wire [22:0] x0;
  wire [23:0] ma;
  wire [22:0] x2;
  wire [7:0] e;
  wire s;
  assign x0=x0reg;
  assign ma=mareg;
  assign x2=x2reg;
  assign e=ereg;
  assign s=sreg;
  
  assign x2wire = tab2(m[22:12]);

  wire [47:0] ax2;
  wire [23:0] ax2_2;
  ///////
  assign ax2 = ma * {1'b1,x2};

  reg [47:0] ax2reg2;
  reg [22:0] x0reg2;
  reg [7:0] ereg2;
  reg sreg2;
 
/////////
  assign ax2_2 = (ax2reg2[47] == 0) ? ax2reg2[46:23] : ax2reg2[47:24];
  
  wire [24:0] x0_2;
  
  assign x0_2 = {1'b1,x0reg2} << 1;
  
  wire [24:0] ans;
  
  assign ans = x0_2 - {1'b0,ax2_2};
  assign y = (ereg2 == 23'b0 || ereg2 == 23'd255) ? {sreg2,31'b0} : ((ereg2 < 8'd253) ? {sreg2,8'd253-ereg2,ans[22:0]} : {s,31'b0});

  always @(posedge clk) begin
    x0reg<=x0wire;
    mareg<=mawire;
    x2reg<=x2wire;
    ereg<=ewire;
    sreg<=swire;

    ax2reg2<=ax2;
    x0reg2<=x0;
    ereg2<=e;
    sreg2<=s;
    
  end

  
endmodule
`default_nettype wire


